module main (input [0:3] Switch,  output [0:3] LED);
       
assign LED = Switch;
 
endmodule
