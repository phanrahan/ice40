// Reading file 'blink.asc'..

module chip (input io_0_8_1, output io_13_9_1);

wire io_0_8_1;
// (0, 0, 'glb_netwk_6')
// (0, 8, 'fabout')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'local_g1_4')
// (0, 8, 'span4_horz_12')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 8, 'sp4_h_r_25')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (2, 8, 'sp4_h_r_36')
// (3, 8, 'sp4_h_l_36')
// (11, 6, 'lutff_global/clk')
// (12, 6, 'lutff_global/clk')
// (12, 7, 'lutff_global/clk')
// (12, 8, 'lutff_global/clk')

reg n2 = 0;
// (10, 5, 'neigh_op_tnr_3')
// (10, 6, 'neigh_op_rgt_3')
// (10, 7, 'neigh_op_bnr_3')
// (11, 5, 'neigh_op_top_3')
// (11, 6, 'local_g0_3')
// (11, 6, 'lutff_3/in_0')
// (11, 6, 'lutff_3/out')
// (11, 7, 'neigh_op_bot_3')
// (12, 5, 'neigh_op_tnl_3')
// (12, 6, 'local_g1_3')
// (12, 6, 'lutff_0/in_2')
// (12, 6, 'lutff_1/in_3')
// (12, 6, 'neigh_op_lft_3')
// (12, 7, 'neigh_op_bnl_3')

reg n3 = 0;
// (11, 5, 'neigh_op_tnr_1')
// (11, 6, 'neigh_op_rgt_1')
// (11, 7, 'neigh_op_bnr_1')
// (12, 5, 'neigh_op_top_1')
// (12, 6, 'local_g3_1')
// (12, 6, 'lutff_1/in_1')
// (12, 6, 'lutff_1/out')
// (12, 7, 'neigh_op_bot_1')
// (13, 5, 'logic_op_tnl_1')
// (13, 6, 'logic_op_lft_1')
// (13, 7, 'logic_op_bnl_1')

reg n4 = 0;
// (11, 5, 'neigh_op_tnr_2')
// (11, 6, 'neigh_op_rgt_2')
// (11, 7, 'neigh_op_bnr_2')
// (12, 5, 'neigh_op_top_2')
// (12, 6, 'local_g3_2')
// (12, 6, 'lutff_2/in_1')
// (12, 6, 'lutff_2/out')
// (12, 7, 'neigh_op_bot_2')
// (13, 5, 'logic_op_tnl_2')
// (13, 6, 'logic_op_lft_2')
// (13, 7, 'logic_op_bnl_2')

reg n5 = 0;
// (11, 5, 'neigh_op_tnr_3')
// (11, 6, 'neigh_op_rgt_3')
// (11, 7, 'neigh_op_bnr_3')
// (12, 5, 'neigh_op_top_3')
// (12, 6, 'local_g0_3')
// (12, 6, 'lutff_3/in_2')
// (12, 6, 'lutff_3/out')
// (12, 7, 'neigh_op_bot_3')
// (13, 5, 'logic_op_tnl_3')
// (13, 6, 'logic_op_lft_3')
// (13, 7, 'logic_op_bnl_3')

reg n6 = 0;
// (11, 5, 'neigh_op_tnr_4')
// (11, 6, 'neigh_op_rgt_4')
// (11, 7, 'neigh_op_bnr_4')
// (12, 5, 'neigh_op_top_4')
// (12, 6, 'local_g0_4')
// (12, 6, 'lutff_4/in_2')
// (12, 6, 'lutff_4/out')
// (12, 7, 'neigh_op_bot_4')
// (13, 5, 'logic_op_tnl_4')
// (13, 6, 'logic_op_lft_4')
// (13, 7, 'logic_op_bnl_4')

reg n7 = 0;
// (11, 5, 'neigh_op_tnr_5')
// (11, 6, 'neigh_op_rgt_5')
// (11, 7, 'neigh_op_bnr_5')
// (12, 5, 'neigh_op_top_5')
// (12, 6, 'local_g1_5')
// (12, 6, 'lutff_5/in_1')
// (12, 6, 'lutff_5/out')
// (12, 7, 'neigh_op_bot_5')
// (13, 5, 'logic_op_tnl_5')
// (13, 6, 'logic_op_lft_5')
// (13, 7, 'logic_op_bnl_5')

reg n8 = 0;
// (11, 5, 'neigh_op_tnr_6')
// (11, 6, 'neigh_op_rgt_6')
// (11, 7, 'neigh_op_bnr_6')
// (12, 5, 'neigh_op_top_6')
// (12, 6, 'local_g1_6')
// (12, 6, 'lutff_6/in_1')
// (12, 6, 'lutff_6/out')
// (12, 7, 'neigh_op_bot_6')
// (13, 5, 'logic_op_tnl_6')
// (13, 6, 'logic_op_lft_6')
// (13, 7, 'logic_op_bnl_6')

reg n9 = 0;
// (11, 5, 'neigh_op_tnr_7')
// (11, 6, 'neigh_op_rgt_7')
// (11, 7, 'neigh_op_bnr_7')
// (12, 5, 'neigh_op_top_7')
// (12, 6, 'local_g3_7')
// (12, 6, 'lutff_7/in_1')
// (12, 6, 'lutff_7/out')
// (12, 7, 'neigh_op_bot_7')
// (13, 5, 'logic_op_tnl_7')
// (13, 6, 'logic_op_lft_7')
// (13, 7, 'logic_op_bnl_7')

reg n10 = 0;
// (11, 6, 'neigh_op_tnr_0')
// (11, 7, 'neigh_op_rgt_0')
// (11, 8, 'neigh_op_bnr_0')
// (12, 6, 'neigh_op_top_0')
// (12, 7, 'local_g3_0')
// (12, 7, 'lutff_0/in_1')
// (12, 7, 'lutff_0/out')
// (12, 8, 'neigh_op_bot_0')
// (13, 6, 'logic_op_tnl_0')
// (13, 7, 'logic_op_lft_0')
// (13, 8, 'logic_op_bnl_0')

reg n11 = 0;
// (11, 6, 'neigh_op_tnr_1')
// (11, 7, 'neigh_op_rgt_1')
// (11, 8, 'neigh_op_bnr_1')
// (12, 6, 'neigh_op_top_1')
// (12, 7, 'local_g0_1')
// (12, 7, 'lutff_1/in_2')
// (12, 7, 'lutff_1/out')
// (12, 8, 'neigh_op_bot_1')
// (13, 6, 'logic_op_tnl_1')
// (13, 7, 'logic_op_lft_1')
// (13, 8, 'logic_op_bnl_1')

reg n12 = 0;
// (11, 6, 'neigh_op_tnr_2')
// (11, 7, 'neigh_op_rgt_2')
// (11, 8, 'neigh_op_bnr_2')
// (12, 6, 'neigh_op_top_2')
// (12, 7, 'local_g0_2')
// (12, 7, 'lutff_2/in_2')
// (12, 7, 'lutff_2/out')
// (12, 8, 'neigh_op_bot_2')
// (13, 6, 'logic_op_tnl_2')
// (13, 7, 'logic_op_lft_2')
// (13, 8, 'logic_op_bnl_2')

reg n13 = 0;
// (11, 6, 'neigh_op_tnr_3')
// (11, 7, 'neigh_op_rgt_3')
// (11, 8, 'neigh_op_bnr_3')
// (12, 6, 'neigh_op_top_3')
// (12, 7, 'local_g0_3')
// (12, 7, 'lutff_3/in_2')
// (12, 7, 'lutff_3/out')
// (12, 8, 'neigh_op_bot_3')
// (13, 6, 'logic_op_tnl_3')
// (13, 7, 'logic_op_lft_3')
// (13, 8, 'logic_op_bnl_3')

reg n14 = 0;
// (11, 6, 'neigh_op_tnr_4')
// (11, 7, 'neigh_op_rgt_4')
// (11, 8, 'neigh_op_bnr_4')
// (12, 6, 'neigh_op_top_4')
// (12, 7, 'local_g2_4')
// (12, 7, 'lutff_4/in_2')
// (12, 7, 'lutff_4/out')
// (12, 8, 'neigh_op_bot_4')
// (13, 6, 'logic_op_tnl_4')
// (13, 7, 'logic_op_lft_4')
// (13, 8, 'logic_op_bnl_4')

reg n15 = 0;
// (11, 6, 'neigh_op_tnr_5')
// (11, 7, 'neigh_op_rgt_5')
// (11, 8, 'neigh_op_bnr_5')
// (12, 6, 'neigh_op_top_5')
// (12, 7, 'local_g2_5')
// (12, 7, 'lutff_5/in_2')
// (12, 7, 'lutff_5/out')
// (12, 8, 'neigh_op_bot_5')
// (13, 6, 'logic_op_tnl_5')
// (13, 7, 'logic_op_lft_5')
// (13, 8, 'logic_op_bnl_5')

reg n16 = 0;
// (11, 6, 'neigh_op_tnr_6')
// (11, 7, 'neigh_op_rgt_6')
// (11, 8, 'neigh_op_bnr_6')
// (12, 6, 'neigh_op_top_6')
// (12, 7, 'local_g0_6')
// (12, 7, 'lutff_6/in_2')
// (12, 7, 'lutff_6/out')
// (12, 8, 'neigh_op_bot_6')
// (13, 6, 'logic_op_tnl_6')
// (13, 7, 'logic_op_lft_6')
// (13, 8, 'logic_op_bnl_6')

reg n17 = 0;
// (11, 6, 'neigh_op_tnr_7')
// (11, 7, 'neigh_op_rgt_7')
// (11, 8, 'neigh_op_bnr_7')
// (12, 6, 'neigh_op_top_7')
// (12, 7, 'local_g1_7')
// (12, 7, 'lutff_7/in_1')
// (12, 7, 'lutff_7/out')
// (12, 8, 'neigh_op_bot_7')
// (13, 6, 'logic_op_tnl_7')
// (13, 7, 'logic_op_lft_7')
// (13, 8, 'logic_op_bnl_7')

reg n18 = 0;
// (11, 7, 'neigh_op_tnr_0')
// (11, 8, 'neigh_op_rgt_0')
// (11, 9, 'neigh_op_bnr_0')
// (12, 7, 'neigh_op_top_0')
// (12, 8, 'local_g2_0')
// (12, 8, 'lutff_0/in_2')
// (12, 8, 'lutff_0/out')
// (12, 9, 'neigh_op_bot_0')
// (13, 7, 'logic_op_tnl_0')
// (13, 8, 'logic_op_lft_0')
// (13, 9, 'logic_op_bnl_0')

reg n19 = 0;
// (11, 7, 'neigh_op_tnr_1')
// (11, 8, 'neigh_op_rgt_1')
// (11, 9, 'neigh_op_bnr_1')
// (12, 7, 'neigh_op_top_1')
// (12, 8, 'local_g3_1')
// (12, 8, 'lutff_1/in_1')
// (12, 8, 'lutff_1/out')
// (12, 9, 'neigh_op_bot_1')
// (13, 7, 'logic_op_tnl_1')
// (13, 8, 'logic_op_lft_1')
// (13, 9, 'logic_op_bnl_1')

reg n20 = 0;
// (11, 7, 'neigh_op_tnr_2')
// (11, 8, 'neigh_op_rgt_2')
// (11, 9, 'neigh_op_bnr_2')
// (12, 7, 'neigh_op_top_2')
// (12, 8, 'local_g3_2')
// (12, 8, 'lutff_2/in_1')
// (12, 8, 'lutff_2/out')
// (12, 9, 'neigh_op_bot_2')
// (13, 7, 'logic_op_tnl_2')
// (13, 8, 'logic_op_lft_2')
// (13, 9, 'logic_op_bnl_2')

reg n21 = 0;
// (11, 7, 'neigh_op_tnr_3')
// (11, 8, 'neigh_op_rgt_3')
// (11, 9, 'neigh_op_bnr_3')
// (12, 7, 'neigh_op_top_3')
// (12, 8, 'local_g1_3')
// (12, 8, 'lutff_3/in_1')
// (12, 8, 'lutff_3/out')
// (12, 9, 'neigh_op_bot_3')
// (13, 7, 'logic_op_tnl_3')
// (13, 8, 'logic_op_lft_3')
// (13, 9, 'logic_op_bnl_3')

reg n22 = 0;
// (11, 7, 'neigh_op_tnr_4')
// (11, 8, 'neigh_op_rgt_4')
// (11, 9, 'neigh_op_bnr_4')
// (12, 7, 'neigh_op_top_4')
// (12, 8, 'local_g1_4')
// (12, 8, 'lutff_4/in_1')
// (12, 8, 'lutff_4/out')
// (12, 9, 'neigh_op_bot_4')
// (13, 7, 'logic_op_tnl_4')
// (13, 8, 'logic_op_lft_4')
// (13, 9, 'logic_op_bnl_4')

reg n23 = 0;
// (11, 7, 'neigh_op_tnr_5')
// (11, 8, 'neigh_op_rgt_5')
// (11, 9, 'neigh_op_bnr_5')
// (12, 7, 'neigh_op_top_5')
// (12, 8, 'local_g2_5')
// (12, 8, 'lutff_5/in_2')
// (12, 8, 'lutff_5/out')
// (12, 9, 'neigh_op_bot_5')
// (13, 7, 'logic_op_tnl_5')
// (13, 8, 'logic_op_lft_5')
// (13, 9, 'logic_op_bnl_5')

reg n24 = 0;
// (11, 7, 'neigh_op_tnr_6')
// (11, 8, 'neigh_op_rgt_6')
// (11, 9, 'neigh_op_bnr_6')
// (12, 7, 'neigh_op_top_6')
// (12, 8, 'local_g1_6')
// (12, 8, 'lutff_6/in_1')
// (12, 8, 'lutff_6/out')
// (12, 9, 'neigh_op_bot_6')
// (13, 7, 'logic_op_tnl_6')
// (13, 8, 'logic_op_lft_6')
// (13, 9, 'logic_op_bnl_6')

reg io_13_9_1 = 0;
// (11, 7, 'neigh_op_tnr_7')
// (11, 8, 'neigh_op_rgt_7')
// (11, 9, 'neigh_op_bnr_7')
// (12, 7, 'neigh_op_top_7')
// (12, 8, 'local_g3_7')
// (12, 8, 'lutff_7/in_1')
// (12, 8, 'lutff_7/out')
// (12, 9, 'neigh_op_bot_7')
// (13, 7, 'logic_op_tnl_7')
// (13, 8, 'logic_op_lft_7')
// (13, 9, 'io_1/D_OUT_0')
// (13, 9, 'io_1/PAD')
// (13, 9, 'local_g0_7')
// (13, 9, 'logic_op_bnl_7')

wire n26;
// (12, 6, 'lutff_1/cout')
// (12, 6, 'lutff_2/in_3')

wire n27;
// (12, 6, 'lutff_2/cout')
// (12, 6, 'lutff_3/in_3')

wire n28;
// (12, 6, 'lutff_3/cout')
// (12, 6, 'lutff_4/in_3')

wire n29;
// (12, 6, 'lutff_4/cout')
// (12, 6, 'lutff_5/in_3')

wire n30;
// (12, 6, 'lutff_5/cout')
// (12, 6, 'lutff_6/in_3')

wire n31;
// (12, 6, 'lutff_6/cout')
// (12, 6, 'lutff_7/in_3')

wire n32;
// (12, 6, 'lutff_7/cout')
// (12, 7, 'carry_in')
// (12, 7, 'carry_in_mux')
// (12, 7, 'lutff_0/in_3')

wire n33;
// (12, 7, 'lutff_0/cout')
// (12, 7, 'lutff_1/in_3')

wire n34;
// (12, 7, 'lutff_1/cout')
// (12, 7, 'lutff_2/in_3')

wire n35;
// (12, 7, 'lutff_2/cout')
// (12, 7, 'lutff_3/in_3')

wire n36;
// (12, 7, 'lutff_3/cout')
// (12, 7, 'lutff_4/in_3')

wire n37;
// (12, 7, 'lutff_4/cout')
// (12, 7, 'lutff_5/in_3')

wire n38;
// (12, 7, 'lutff_5/cout')
// (12, 7, 'lutff_6/in_3')

wire n39;
// (12, 7, 'lutff_6/cout')
// (12, 7, 'lutff_7/in_3')

wire n40;
// (12, 7, 'lutff_7/cout')
// (12, 8, 'carry_in')
// (12, 8, 'carry_in_mux')
// (12, 8, 'lutff_0/in_3')

wire n41;
// (12, 8, 'lutff_0/cout')
// (12, 8, 'lutff_1/in_3')

wire n42;
// (12, 8, 'lutff_1/cout')
// (12, 8, 'lutff_2/in_3')

wire n43;
// (12, 8, 'lutff_2/cout')
// (12, 8, 'lutff_3/in_3')

wire n44;
// (12, 8, 'lutff_3/cout')
// (12, 8, 'lutff_4/in_3')

wire n45;
// (12, 8, 'lutff_4/cout')
// (12, 8, 'lutff_5/in_3')

wire n46;
// (12, 8, 'lutff_5/cout')
// (12, 8, 'lutff_6/in_3')

wire n47;
// (12, 8, 'lutff_6/cout')
// (12, 8, 'lutff_7/in_3')

wire n48;
// (12, 6, 'lutff_0/cout')

wire n49;
// (12, 6, 'lutff_2/lout')

wire n50;
// (12, 7, 'lutff_1/lout')

wire n51;
// (12, 7, 'lutff_7/lout')

wire n52;
// (12, 6, 'lutff_5/lout')

wire n53;
// (12, 8, 'lutff_2/lout')

wire n54;
// (12, 7, 'lutff_4/lout')

wire n55;
// (11, 6, 'lutff_3/lout')

wire n56;
// (12, 8, 'lutff_5/lout')

wire n57;
// (12, 7, 'lutff_0/lout')

wire n58;
// (12, 7, 'lutff_3/lout')

wire n59;
// (12, 6, 'lutff_1/lout')

wire n60;
// (12, 6, 'lutff_7/lout')

wire n61;
// (12, 8, 'lutff_4/lout')

wire n62;
// (12, 7, 'lutff_6/lout')

wire n63;
// (12, 6, 'lutff_4/lout')

wire n64;
// (12, 8, 'lutff_1/lout')

wire n65;
// (12, 8, 'lutff_7/lout')

wire n66;
// (12, 6, 'lutff_0/out')

wire n67;
// (12, 6, 'lutff_0/lout')

wire n68;
// (12, 6, 'carry_in_mux')

// Carry-In for (12 6)
assign n68 = 1;

wire n69;
// (12, 7, 'lutff_5/lout')

wire n70;
// (12, 6, 'lutff_3/lout')

wire n71;
// (12, 8, 'lutff_0/lout')

wire n72;
// (12, 7, 'lutff_2/lout')

wire n73;
// (12, 6, 'lutff_6/lout')

wire n74;
// (12, 8, 'lutff_3/lout')

wire n75;
// (12, 8, 'lutff_6/lout')

assign n67 = /* LUT   12  6  0 */ 1'b0;
assign n49 = /* LUT   12  6  2 */ (n26 ? !n4 : n4);
assign n50 = /* LUT   12  7  1 */ (n33 ? !n11 : n11);
assign n51 = /* LUT   12  7  7 */ (n39 ? !n17 : n17);
assign n52 = /* LUT   12  6  5 */ (n29 ? !n7 : n7);
assign n53 = /* LUT   12  8  2 */ (n42 ? !n20 : n20);
assign n54 = /* LUT   12  7  4 */ (n36 ? !n14 : n14);
assign n55 = /* LUT   11  6  3 */ !n2;
assign n56 = /* LUT   12  8  5 */ (n45 ? !n23 : n23);
assign n57 = /* LUT   12  7  0 */ (n32 ? !n10 : n10);
assign n58 = /* LUT   12  7  3 */ (n35 ? !n13 : n13);
assign n59 = /* LUT   12  6  1 */ (n2 ? !n3 : n3);
assign n60 = /* LUT   12  6  7 */ (n31 ? !n9 : n9);
assign n61 = /* LUT   12  8  4 */ (n44 ? !n22 : n22);
assign n62 = /* LUT   12  7  6 */ (n38 ? !n16 : n16);
assign n63 = /* LUT   12  6  4 */ (n28 ? !n6 : n6);
assign n64 = /* LUT   12  8  1 */ (n41 ? !n19 : n19);
assign n65 = /* LUT   12  8  7 */ (n47 ? !io_13_9_1 : io_13_9_1);
assign n69 = /* LUT   12  7  5 */ (n37 ? !n15 : n15);
assign n70 = /* LUT   12  6  3 */ (n27 ? !n5 : n5);
assign n71 = /* LUT   12  8  0 */ (n40 ? !n18 : n18);
assign n72 = /* LUT   12  7  2 */ (n34 ? !n12 : n12);
assign n73 = /* LUT   12  6  6 */ (n30 ? !n8 : n8);
assign n74 = /* LUT   12  8  3 */ (n43 ? !n21 : n21);
assign n75 = /* LUT   12  8  6 */ (n46 ? !n24 : n24);
assign n27 = /* CARRY 12  6  2 */ (n4 & 1'b0) | ((n4 | 1'b0) & n26);
assign n34 = /* CARRY 12  7  1 */ (1'b0 & n11) | ((1'b0 | n11) & n33);
assign n40 = /* CARRY 12  7  7 */ (n17 & 1'b0) | ((n17 | 1'b0) & n39);
assign n30 = /* CARRY 12  6  5 */ (n7 & 1'b0) | ((n7 | 1'b0) & n29);
assign n43 = /* CARRY 12  8  2 */ (n20 & 1'b0) | ((n20 | 1'b0) & n42);
assign n37 = /* CARRY 12  7  4 */ (1'b0 & n14) | ((1'b0 | n14) & n36);
assign n46 = /* CARRY 12  8  5 */ (1'b0 & n23) | ((1'b0 | n23) & n45);
assign n33 = /* CARRY 12  7  0 */ (n10 & 1'b0) | ((n10 | 1'b0) & n32);
assign n36 = /* CARRY 12  7  3 */ (1'b0 & n13) | ((1'b0 | n13) & n35);
assign n26 = /* CARRY 12  6  1 */ (n3 & 1'b0) | ((n3 | 1'b0) & n48);
assign n32 = /* CARRY 12  6  7 */ (n9 & 1'b0) | ((n9 | 1'b0) & n31);
assign n45 = /* CARRY 12  8  4 */ (n22 & 1'b0) | ((n22 | 1'b0) & n44);
assign n39 = /* CARRY 12  7  6 */ (1'b0 & n16) | ((1'b0 | n16) & n38);
assign n29 = /* CARRY 12  6  4 */ (1'b0 & n6) | ((1'b0 | n6) & n28);
assign n42 = /* CARRY 12  8  1 */ (n19 & 1'b0) | ((n19 | 1'b0) & n41);
assign n48 = /* CARRY 12  6  0 */ (1'b0 & n2) | ((1'b0 | n2) & n68);
assign n38 = /* CARRY 12  7  5 */ (1'b0 & n15) | ((1'b0 | n15) & n37);
assign n28 = /* CARRY 12  6  3 */ (1'b0 & n5) | ((1'b0 | n5) & n27);
assign n41 = /* CARRY 12  8  0 */ (1'b0 & n18) | ((1'b0 | n18) & n40);
assign n35 = /* CARRY 12  7  2 */ (1'b0 & n12) | ((1'b0 | n12) & n34);
assign n31 = /* CARRY 12  6  6 */ (n8 & 1'b0) | ((n8 | 1'b0) & n30);
assign n44 = /* CARRY 12  8  3 */ (n21 & 1'b0) | ((n21 | 1'b0) & n43);
assign n47 = /* CARRY 12  8  6 */ (n24 & 1'b0) | ((n24 | 1'b0) & n46);
/* FF 12  6  2 */ always @(posedge io_0_8_1) if (1'b1) n4 <= 1'b0 ? 1'b0 : n49;
/* FF 12  7  1 */ always @(posedge io_0_8_1) if (1'b1) n11 <= 1'b0 ? 1'b0 : n50;
/* FF 12  7  7 */ always @(posedge io_0_8_1) if (1'b1) n17 <= 1'b0 ? 1'b0 : n51;
/* FF 12  6  5 */ always @(posedge io_0_8_1) if (1'b1) n7 <= 1'b0 ? 1'b0 : n52;
/* FF 12  8  2 */ always @(posedge io_0_8_1) if (1'b1) n20 <= 1'b0 ? 1'b0 : n53;
/* FF 12  7  4 */ always @(posedge io_0_8_1) if (1'b1) n14 <= 1'b0 ? 1'b0 : n54;
/* FF 11  6  3 */ always @(posedge io_0_8_1) if (1'b1) n2 <= 1'b0 ? 1'b0 : n55;
/* FF 12  8  5 */ always @(posedge io_0_8_1) if (1'b1) n23 <= 1'b0 ? 1'b0 : n56;
/* FF 12  7  0 */ always @(posedge io_0_8_1) if (1'b1) n10 <= 1'b0 ? 1'b0 : n57;
/* FF 12  7  3 */ always @(posedge io_0_8_1) if (1'b1) n13 <= 1'b0 ? 1'b0 : n58;
/* FF 12  6  1 */ always @(posedge io_0_8_1) if (1'b1) n3 <= 1'b0 ? 1'b0 : n59;
/* FF 12  6  7 */ always @(posedge io_0_8_1) if (1'b1) n9 <= 1'b0 ? 1'b0 : n60;
/* FF 12  8  4 */ always @(posedge io_0_8_1) if (1'b1) n22 <= 1'b0 ? 1'b0 : n61;
/* FF 12  7  6 */ always @(posedge io_0_8_1) if (1'b1) n16 <= 1'b0 ? 1'b0 : n62;
/* FF 12  6  4 */ always @(posedge io_0_8_1) if (1'b1) n6 <= 1'b0 ? 1'b0 : n63;
/* FF 12  8  1 */ always @(posedge io_0_8_1) if (1'b1) n19 <= 1'b0 ? 1'b0 : n64;
/* FF 12  8  7 */ always @(posedge io_0_8_1) if (1'b1) io_13_9_1 <= 1'b0 ? 1'b0 : n65;
/* FF 12  6  0 */ assign n66 = n67;
/* FF 12  7  5 */ always @(posedge io_0_8_1) if (1'b1) n15 <= 1'b0 ? 1'b0 : n69;
/* FF 12  6  3 */ always @(posedge io_0_8_1) if (1'b1) n5 <= 1'b0 ? 1'b0 : n70;
/* FF 12  8  0 */ always @(posedge io_0_8_1) if (1'b1) n18 <= 1'b0 ? 1'b0 : n71;
/* FF 12  7  2 */ always @(posedge io_0_8_1) if (1'b1) n12 <= 1'b0 ? 1'b0 : n72;
/* FF 12  6  6 */ always @(posedge io_0_8_1) if (1'b1) n8 <= 1'b0 ? 1'b0 : n73;
/* FF 12  8  3 */ always @(posedge io_0_8_1) if (1'b1) n21 <= 1'b0 ? 1'b0 : n74;
/* FF 12  8  6 */ always @(posedge io_0_8_1) if (1'b1) n24 <= 1'b0 ? 1'b0 : n75;

endmodule

