// Reading file 'vga.asc'..

module chip (input io_0_8_1, output io_2_0_0, output io_3_0_0, output io_3_0_1, output io_4_0_0, output io_6_0_0, output io_6_0_1, output io_7_0_1, output io_9_0_1, output io_10_0_0, output io_10_0_1, output io_2_0_1);

wire io_0_8_1;
// (0, 0, 'glb_netwk_6')
// (0, 8, 'fabout')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'local_g1_4')
// (0, 8, 'span4_horz_4')
// (1, 2, 'lutff_global/clk')
// (1, 4, 'lutff_global/clk')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 8, 'sp4_h_r_17')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (2, 3, 'lutff_global/clk')
// (2, 4, 'lutff_global/clk')
// (2, 8, 'sp4_h_r_28')
// (3, 8, 'sp4_h_r_41')
// (4, 3, 'lutff_global/clk')
// (4, 4, 'lutff_global/clk')
// (4, 5, 'lutff_global/clk')
// (4, 8, 'sp4_h_l_41')
// (5, 5, 'lutff_global/clk')
// (7, 4, 'lutff_global/clk')

reg io_2_0_0 = 0;
// (0, 1, 'logic_op_tnr_4')
// (0, 2, 'logic_op_rgt_4')
// (0, 3, 'logic_op_bnr_4')
// (1, 1, 'neigh_op_top_4')
// (1, 1, 'sp4_r_v_b_20')
// (1, 2, 'lutff_4/out')
// (1, 2, 'sp4_r_v_b_9')
// (1, 3, 'neigh_op_bot_4')
// (2, 0, 'io_0/D_OUT_0')
// (2, 0, 'io_0/PAD')
// (2, 0, 'local_g0_4')
// (2, 0, 'span4_vert_20')
// (2, 1, 'neigh_op_tnl_4')
// (2, 1, 'sp4_v_b_20')
// (2, 2, 'neigh_op_lft_4')
// (2, 2, 'sp4_v_b_9')
// (2, 3, 'neigh_op_bnl_4')

wire n3;
// (0, 2, 'logic_op_tnr_1')
// (0, 3, 'logic_op_rgt_1')
// (0, 4, 'logic_op_bnr_1')
// (1, 0, 'span4_vert_26')
// (1, 1, 'local_g3_2')
// (1, 1, 'lutff_1/in_2')
// (1, 1, 'sp4_v_b_26')
// (1, 2, 'neigh_op_top_1')
// (1, 2, 'sp4_v_b_15')
// (1, 3, 'local_g3_1')
// (1, 3, 'lutff_1/in_1')
// (1, 3, 'lutff_1/out')
// (1, 3, 'sp4_v_b_2')
// (1, 4, 'neigh_op_bot_1')
// (2, 2, 'neigh_op_tnl_1')
// (2, 3, 'neigh_op_lft_1')
// (2, 4, 'neigh_op_bnl_1')

wire n4;
// (0, 2, 'logic_op_tnr_2')
// (0, 3, 'logic_op_rgt_2')
// (0, 4, 'logic_op_bnr_2')
// (1, 0, 'span4_vert_28')
// (1, 1, 'local_g2_4')
// (1, 1, 'lutff_2/in_2')
// (1, 1, 'sp4_v_b_28')
// (1, 2, 'neigh_op_top_2')
// (1, 2, 'sp4_v_b_17')
// (1, 3, 'local_g2_2')
// (1, 3, 'lutff_2/in_2')
// (1, 3, 'lutff_2/out')
// (1, 3, 'sp4_v_b_4')
// (1, 4, 'neigh_op_bot_2')
// (2, 2, 'neigh_op_tnl_2')
// (2, 3, 'neigh_op_lft_2')
// (2, 4, 'neigh_op_bnl_2')

wire n5;
// (0, 2, 'logic_op_tnr_3')
// (0, 3, 'logic_op_rgt_3')
// (0, 4, 'logic_op_bnr_3')
// (1, 0, 'span4_vert_30')
// (1, 1, 'local_g2_6')
// (1, 1, 'lutff_3/in_1')
// (1, 1, 'sp4_v_b_30')
// (1, 2, 'neigh_op_top_3')
// (1, 2, 'sp4_v_b_19')
// (1, 3, 'local_g1_3')
// (1, 3, 'lutff_3/in_1')
// (1, 3, 'lutff_3/out')
// (1, 3, 'sp4_v_b_6')
// (1, 4, 'neigh_op_bot_3')
// (2, 2, 'neigh_op_tnl_3')
// (2, 3, 'neigh_op_lft_3')
// (2, 4, 'neigh_op_bnl_3')

wire n6;
// (0, 2, 'logic_op_tnr_4')
// (0, 3, 'logic_op_rgt_4')
// (0, 4, 'logic_op_bnr_4')
// (1, 0, 'span4_vert_32')
// (1, 1, 'local_g3_0')
// (1, 1, 'lutff_4/in_1')
// (1, 1, 'sp4_v_b_32')
// (1, 2, 'neigh_op_top_4')
// (1, 2, 'sp4_v_b_21')
// (1, 3, 'local_g1_4')
// (1, 3, 'lutff_4/in_1')
// (1, 3, 'lutff_4/out')
// (1, 3, 'sp4_v_b_8')
// (1, 4, 'neigh_op_bot_4')
// (2, 2, 'neigh_op_tnl_4')
// (2, 3, 'neigh_op_lft_4')
// (2, 4, 'neigh_op_bnl_4')

wire n7;
// (0, 2, 'logic_op_tnr_5')
// (0, 3, 'logic_op_rgt_5')
// (0, 4, 'logic_op_bnr_5')
// (1, 0, 'span4_vert_34')
// (1, 1, 'local_g2_2')
// (1, 1, 'lutff_5/in_1')
// (1, 1, 'sp4_v_b_34')
// (1, 1, 'sp4_v_t_39')
// (1, 2, 'neigh_op_top_5')
// (1, 2, 'sp4_v_b_23')
// (1, 2, 'sp4_v_b_39')
// (1, 3, 'local_g0_5')
// (1, 3, 'lutff_5/in_2')
// (1, 3, 'lutff_5/out')
// (1, 3, 'sp4_v_b_10')
// (1, 3, 'sp4_v_b_26')
// (1, 4, 'neigh_op_bot_5')
// (1, 4, 'sp4_v_b_15')
// (1, 5, 'local_g1_2')
// (1, 5, 'lutff_0/in_1')
// (1, 5, 'sp4_v_b_2')
// (2, 2, 'neigh_op_tnl_5')
// (2, 3, 'neigh_op_lft_5')
// (2, 4, 'neigh_op_bnl_5')

wire n8;
// (0, 2, 'logic_op_tnr_6')
// (0, 3, 'logic_op_rgt_6')
// (0, 4, 'logic_op_bnr_6')
// (1, 0, 'span4_vert_36')
// (1, 1, 'local_g3_4')
// (1, 1, 'lutff_6/in_1')
// (1, 1, 'sp4_v_b_36')
// (1, 2, 'neigh_op_top_6')
// (1, 2, 'sp4_v_b_25')
// (1, 3, 'local_g2_6')
// (1, 3, 'lutff_6/in_2')
// (1, 3, 'lutff_6/out')
// (1, 3, 'sp4_r_v_b_45')
// (1, 3, 'sp4_v_b_12')
// (1, 4, 'neigh_op_bot_6')
// (1, 4, 'sp4_r_v_b_32')
// (1, 4, 'sp4_v_b_1')
// (1, 5, 'local_g3_5')
// (1, 5, 'lutff_1/in_1')
// (1, 5, 'sp4_r_v_b_21')
// (1, 6, 'sp4_r_v_b_8')
// (2, 2, 'neigh_op_tnl_6')
// (2, 2, 'sp4_v_t_45')
// (2, 3, 'neigh_op_lft_6')
// (2, 3, 'sp4_v_b_45')
// (2, 4, 'neigh_op_bnl_6')
// (2, 4, 'sp4_v_b_32')
// (2, 5, 'sp4_v_b_21')
// (2, 6, 'sp4_v_b_8')

wire n9;
// (0, 2, 'logic_op_tnr_7')
// (0, 3, 'logic_op_rgt_7')
// (0, 4, 'logic_op_bnr_7')
// (1, 0, 'span4_vert_38')
// (1, 1, 'local_g3_6')
// (1, 1, 'lutff_7/in_2')
// (1, 1, 'sp4_v_b_38')
// (1, 2, 'neigh_op_top_7')
// (1, 2, 'sp4_v_b_27')
// (1, 2, 'sp4_v_t_46')
// (1, 3, 'local_g1_7')
// (1, 3, 'lutff_7/in_1')
// (1, 3, 'lutff_7/out')
// (1, 3, 'sp4_v_b_14')
// (1, 3, 'sp4_v_b_46')
// (1, 4, 'neigh_op_bot_7')
// (1, 4, 'sp4_v_b_3')
// (1, 4, 'sp4_v_b_35')
// (1, 5, 'local_g0_6')
// (1, 5, 'lutff_2/in_2')
// (1, 5, 'sp4_v_b_22')
// (1, 6, 'sp4_v_b_11')
// (2, 2, 'neigh_op_tnl_7')
// (2, 3, 'neigh_op_lft_7')
// (2, 4, 'neigh_op_bnl_7')

wire n10;
// (0, 3, 'logic_op_tnr_0')
// (0, 4, 'logic_op_rgt_0')
// (0, 5, 'logic_op_bnr_0')
// (1, 0, 'span4_vert_37')
// (1, 1, 'sp4_v_b_37')
// (1, 2, 'local_g2_0')
// (1, 2, 'lutff_0/in_2')
// (1, 2, 'sp4_v_b_24')
// (1, 3, 'neigh_op_top_0')
// (1, 3, 'sp4_v_b_13')
// (1, 4, 'local_g0_0')
// (1, 4, 'lutff_0/in_2')
// (1, 4, 'lutff_0/out')
// (1, 4, 'sp4_v_b_0')
// (1, 5, 'local_g1_0')
// (1, 5, 'lutff_3/in_2')
// (1, 5, 'neigh_op_bot_0')
// (2, 3, 'neigh_op_tnl_0')
// (2, 4, 'neigh_op_lft_0')
// (2, 5, 'neigh_op_bnl_0')

wire n11;
// (0, 3, 'logic_op_tnr_1')
// (0, 4, 'logic_op_rgt_1')
// (0, 4, 'span4_horz_23')
// (0, 5, 'logic_op_bnr_1')
// (1, 0, 'span12_vert_9')
// (1, 0, 'span4_vert_39')
// (1, 1, 'local_g3_1')
// (1, 1, 'lutff_6/in_2')
// (1, 1, 'lutff_7/in_1')
// (1, 1, 'sp12_v_b_9')
// (1, 1, 'sp4_v_b_39')
// (1, 2, 'local_g3_2')
// (1, 2, 'lutff_1/in_2')
// (1, 2, 'sp12_v_b_6')
// (1, 2, 'sp4_v_b_26')
// (1, 3, 'local_g0_1')
// (1, 3, 'lutff_7/in_2')
// (1, 3, 'neigh_op_top_1')
// (1, 3, 'sp12_v_b_5')
// (1, 3, 'sp4_v_b_15')
// (1, 4, 'local_g1_1')
// (1, 4, 'lutff_1/in_1')
// (1, 4, 'lutff_1/out')
// (1, 4, 'sp12_v_b_2')
// (1, 4, 'sp4_h_r_2')
// (1, 4, 'sp4_h_r_34')
// (1, 4, 'sp4_v_b_2')
// (1, 5, 'local_g0_1')
// (1, 5, 'local_g1_1')
// (1, 5, 'lutff_3/in_1')
// (1, 5, 'lutff_4/in_1')
// (1, 5, 'neigh_op_bot_1')
// (1, 5, 'sp12_v_b_1')
// (2, 3, 'neigh_op_tnl_1')
// (2, 4, 'neigh_op_lft_1')
// (2, 4, 'sp4_h_r_15')
// (2, 4, 'sp4_h_r_47')
// (2, 5, 'neigh_op_bnl_1')
// (3, 4, 'sp4_h_l_47')
// (3, 4, 'sp4_h_r_1')
// (3, 4, 'sp4_h_r_26')
// (4, 1, 'sp4_r_v_b_45')
// (4, 2, 'sp4_r_v_b_32')
// (4, 3, 'sp4_r_v_b_21')
// (4, 4, 'sp4_h_r_12')
// (4, 4, 'sp4_h_r_39')
// (4, 4, 'sp4_r_v_b_8')
// (5, 0, 'span4_vert_45')
// (5, 1, 'sp4_v_b_45')
// (5, 2, 'sp4_v_b_32')
// (5, 3, 'local_g0_5')
// (5, 3, 'local_g1_5')
// (5, 3, 'lutff_2/in_1')
// (5, 3, 'lutff_3/in_1')
// (5, 3, 'sp4_v_b_21')
// (5, 4, 'local_g3_1')
// (5, 4, 'lutff_1/in_1')
// (5, 4, 'sp4_h_l_39')
// (5, 4, 'sp4_h_r_25')
// (5, 4, 'sp4_h_r_5')
// (5, 4, 'sp4_v_b_8')
// (6, 1, 'sp4_r_v_b_36')
// (6, 2, 'sp4_r_v_b_25')
// (6, 3, 'local_g2_4')
// (6, 3, 'lutff_5/in_1')
// (6, 3, 'lutff_6/in_2')
// (6, 3, 'lutff_7/in_1')
// (6, 3, 'sp4_r_v_b_12')
// (6, 4, 'local_g1_0')
// (6, 4, 'lutff_0/in_1')
// (6, 4, 'sp4_h_r_16')
// (6, 4, 'sp4_h_r_36')
// (6, 4, 'sp4_r_v_b_1')
// (7, 0, 'span4_vert_36')
// (7, 1, 'sp4_v_b_36')
// (7, 2, 'sp4_v_b_25')
// (7, 3, 'local_g1_4')
// (7, 3, 'lutff_1/in_2')
// (7, 3, 'lutff_7/in_2')
// (7, 3, 'sp4_v_b_12')
// (7, 4, 'sp4_h_l_36')
// (7, 4, 'sp4_h_r_29')
// (7, 4, 'sp4_v_b_1')
// (8, 4, 'sp4_h_r_40')
// (9, 4, 'sp4_h_l_40')

wire n12;
// (0, 3, 'logic_op_tnr_2')
// (0, 4, 'logic_op_rgt_2')
// (0, 5, 'logic_op_bnr_2')
// (1, 0, 'span4_vert_41')
// (1, 1, 'sp4_v_b_41')
// (1, 2, 'local_g3_4')
// (1, 2, 'lutff_2/in_1')
// (1, 2, 'sp4_v_b_28')
// (1, 3, 'neigh_op_top_2')
// (1, 3, 'sp4_v_b_17')
// (1, 4, 'local_g0_2')
// (1, 4, 'lutff_2/in_2')
// (1, 4, 'lutff_2/out')
// (1, 4, 'sp4_v_b_4')
// (1, 5, 'local_g0_2')
// (1, 5, 'lutff_5/in_1')
// (1, 5, 'neigh_op_bot_2')
// (2, 3, 'neigh_op_tnl_2')
// (2, 4, 'neigh_op_lft_2')
// (2, 5, 'neigh_op_bnl_2')

wire n13;
// (0, 3, 'logic_op_tnr_3')
// (0, 4, 'logic_op_rgt_3')
// (0, 5, 'logic_op_bnr_3')
// (1, 0, 'span4_vert_43')
// (1, 1, 'sp4_v_b_43')
// (1, 2, 'local_g3_6')
// (1, 2, 'lutff_3/in_2')
// (1, 2, 'sp4_v_b_30')
// (1, 3, 'neigh_op_top_3')
// (1, 3, 'sp4_v_b_19')
// (1, 4, 'local_g2_3')
// (1, 4, 'lutff_3/in_2')
// (1, 4, 'lutff_3/out')
// (1, 4, 'sp4_v_b_6')
// (1, 5, 'local_g1_3')
// (1, 5, 'lutff_6/in_2')
// (1, 5, 'neigh_op_bot_3')
// (2, 3, 'neigh_op_tnl_3')
// (2, 4, 'neigh_op_lft_3')
// (2, 5, 'neigh_op_bnl_3')

wire n14;
// (0, 3, 'logic_op_tnr_4')
// (0, 4, 'logic_op_rgt_4')
// (0, 5, 'logic_op_bnr_4')
// (1, 3, 'neigh_op_top_4')
// (1, 4, 'lutff_4/out')
// (1, 4, 'sp4_h_r_8')
// (1, 5, 'neigh_op_bot_4')
// (2, 3, 'neigh_op_tnl_4')
// (2, 4, 'neigh_op_lft_4')
// (2, 4, 'sp4_h_r_21')
// (2, 5, 'neigh_op_bnl_4')
// (3, 4, 'sp4_h_r_32')
// (4, 4, 'sp4_h_r_45')
// (5, 4, 'sp4_h_l_45')
// (5, 4, 'sp4_h_r_11')
// (6, 4, 'local_g0_6')
// (6, 4, 'lutff_4/in_0')
// (6, 4, 'sp4_h_r_22')
// (7, 4, 'sp4_h_r_35')
// (8, 4, 'sp4_h_r_46')
// (9, 4, 'sp4_h_l_46')

wire n15;
// (0, 3, 'logic_op_tnr_5')
// (0, 4, 'logic_op_rgt_5')
// (0, 5, 'logic_op_bnr_5')
// (1, 0, 'span4_vert_47')
// (1, 1, 'local_g3_7')
// (1, 1, 'lutff_0/in_2')
// (1, 1, 'sp4_v_b_47')
// (1, 2, 'sp4_v_b_34')
// (1, 3, 'local_g1_5')
// (1, 3, 'lutff_0/in_2')
// (1, 3, 'neigh_op_top_5')
// (1, 3, 'sp4_v_b_23')
// (1, 4, 'local_g2_5')
// (1, 4, 'lutff_5/out')
// (1, 4, 'lutff_6/in_3')
// (1, 4, 'sp4_v_b_10')
// (1, 5, 'neigh_op_bot_5')
// (2, 3, 'neigh_op_tnl_5')
// (2, 4, 'neigh_op_lft_5')
// (2, 5, 'neigh_op_bnl_5')

reg n16 = 0;
// (0, 3, 'logic_op_tnr_6')
// (0, 4, 'logic_op_rgt_6')
// (0, 5, 'logic_op_bnr_6')
// (1, 3, 'neigh_op_top_6')
// (1, 4, 'local_g0_6')
// (1, 4, 'lutff_5/in_3')
// (1, 4, 'lutff_6/out')
// (1, 4, 'lutff_7/in_3')
// (1, 5, 'neigh_op_bot_6')
// (2, 3, 'local_g2_6')
// (2, 3, 'lutff_0/in_2')
// (2, 3, 'neigh_op_tnl_6')
// (2, 4, 'local_g0_6')
// (2, 4, 'lutff_4/in_0')
// (2, 4, 'lutff_7/in_3')
// (2, 4, 'neigh_op_lft_6')
// (2, 5, 'neigh_op_bnl_6')

wire n17;
// (0, 3, 'logic_op_tnr_7')
// (0, 4, 'logic_op_rgt_7')
// (0, 5, 'logic_op_bnr_7')
// (1, 3, 'neigh_op_top_7')
// (1, 4, 'lutff_7/out')
// (1, 5, 'local_g1_7')
// (1, 5, 'lutff_7/in_1')
// (1, 5, 'neigh_op_bot_7')
// (2, 3, 'neigh_op_tnl_7')
// (2, 4, 'neigh_op_lft_7')
// (2, 5, 'neigh_op_bnl_7')

wire n18;
// (0, 4, 'logic_op_tnr_4')
// (0, 5, 'logic_op_rgt_4')
// (0, 6, 'logic_op_bnr_4')
// (1, 1, 'sp4_v_t_45')
// (1, 2, 'local_g3_5')
// (1, 2, 'lutff_1/in_1')
// (1, 2, 'sp4_v_b_45')
// (1, 3, 'sp4_v_b_32')
// (1, 4, 'local_g1_4')
// (1, 4, 'lutff_1/in_2')
// (1, 4, 'neigh_op_top_4')
// (1, 4, 'sp4_v_b_21')
// (1, 5, 'local_g2_4')
// (1, 5, 'lutff_4/in_2')
// (1, 5, 'lutff_4/out')
// (1, 5, 'sp4_v_b_8')
// (1, 6, 'neigh_op_bot_4')
// (2, 4, 'neigh_op_tnl_4')
// (2, 5, 'neigh_op_lft_4')
// (2, 6, 'neigh_op_bnl_4')

wire n19;
// (0, 4, 'logic_op_tnr_7')
// (0, 5, 'logic_op_rgt_7')
// (0, 5, 'span4_horz_3')
// (0, 5, 'span4_horz_35')
// (0, 6, 'logic_op_bnr_7')
// (1, 2, 'sp4_r_v_b_40')
// (1, 3, 'sp4_r_v_b_29')
// (1, 4, 'local_g0_4')
// (1, 4, 'lutff_global/s_r')
// (1, 4, 'neigh_op_top_7')
// (1, 4, 'sp4_h_r_4')
// (1, 4, 'sp4_r_v_b_16')
// (1, 4, 'sp4_v_t_46')
// (1, 5, 'lutff_7/out')
// (1, 5, 'sp4_h_r_14')
// (1, 5, 'sp4_h_r_46')
// (1, 5, 'sp4_r_v_b_47')
// (1, 5, 'sp4_r_v_b_5')
// (1, 5, 'sp4_v_b_46')
// (1, 6, 'neigh_op_bot_7')
// (1, 6, 'sp4_r_v_b_34')
// (1, 6, 'sp4_v_b_35')
// (1, 7, 'sp4_r_v_b_23')
// (1, 7, 'sp4_v_b_22')
// (1, 8, 'sp4_r_v_b_10')
// (1, 8, 'sp4_v_b_11')
// (2, 1, 'sp4_v_t_40')
// (2, 2, 'sp4_v_b_40')
// (2, 3, 'local_g3_5')
// (2, 3, 'lutff_global/s_r')
// (2, 3, 'sp4_v_b_29')
// (2, 4, 'neigh_op_tnl_7')
// (2, 4, 'sp4_h_r_10')
// (2, 4, 'sp4_h_r_17')
// (2, 4, 'sp4_v_b_16')
// (2, 4, 'sp4_v_t_47')
// (2, 5, 'local_g1_7')
// (2, 5, 'lutff_5/in_1')
// (2, 5, 'neigh_op_lft_7')
// (2, 5, 'sp4_h_l_46')
// (2, 5, 'sp4_h_r_27')
// (2, 5, 'sp4_v_b_47')
// (2, 5, 'sp4_v_b_5')
// (2, 6, 'neigh_op_bnl_7')
// (2, 6, 'sp4_v_b_34')
// (2, 7, 'sp4_v_b_23')
// (2, 8, 'sp4_v_b_10')
// (3, 2, 'sp4_r_v_b_38')
// (3, 3, 'sp4_r_v_b_27')
// (3, 4, 'sp4_h_r_23')
// (3, 4, 'sp4_h_r_28')
// (3, 4, 'sp4_r_v_b_14')
// (3, 5, 'sp4_h_r_38')
// (3, 5, 'sp4_r_v_b_3')
// (4, 1, 'sp4_v_t_38')
// (4, 2, 'sp4_v_b_38')
// (4, 3, 'local_g3_3')
// (4, 3, 'lutff_global/cen')
// (4, 3, 'sp4_v_b_27')
// (4, 4, 'local_g2_2')
// (4, 4, 'lutff_global/cen')
// (4, 4, 'sp4_h_r_34')
// (4, 4, 'sp4_h_r_41')
// (4, 4, 'sp4_v_b_14')
// (4, 5, 'sp4_h_l_38')
// (4, 5, 'sp4_h_r_6')
// (4, 5, 'sp4_v_b_3')
// (5, 4, 'sp4_h_l_41')
// (5, 4, 'sp4_h_r_47')
// (5, 5, 'local_g1_3')
// (5, 5, 'lutff_global/cen')
// (5, 5, 'sp4_h_r_19')
// (6, 4, 'sp4_h_l_47')
// (6, 5, 'sp4_h_r_30')
// (7, 5, 'sp4_h_r_43')
// (8, 5, 'sp4_h_l_43')

reg io_3_0_0 = 0;
assign io_3_0_1 = io_3_0_0;
assign io_4_0_0 = io_3_0_0;
assign io_6_0_0 = io_3_0_0;
assign io_6_0_1 = io_3_0_0;
assign io_7_0_1 = io_3_0_0;
assign io_9_0_1 = io_3_0_0;
assign io_10_0_0 = io_3_0_0;
assign io_10_0_1 = io_3_0_0;
// (0, 5, 'span12_horz_10')
// (1, 0, 'span4_horz_r_1')
// (1, 5, 'sp12_h_r_13')
// (2, 0, 'span4_horz_r_5')
// (2, 5, 'sp12_h_r_14')
// (3, 0, 'io_0/D_OUT_0')
// (3, 0, 'io_0/PAD')
// (3, 0, 'io_1/D_OUT_0')
// (3, 0, 'io_1/PAD')
// (3, 0, 'local_g0_1')
// (3, 0, 'local_g1_1')
// (3, 0, 'span4_horz_r_9')
// (3, 1, 'sp4_r_v_b_6')
// (3, 2, 'sp4_r_v_b_47')
// (3, 3, 'sp4_r_v_b_34')
// (3, 4, 'neigh_op_tnr_5')
// (3, 4, 'sp4_r_v_b_23')
// (3, 5, 'neigh_op_rgt_5')
// (3, 5, 'sp12_h_r_17')
// (3, 5, 'sp4_r_v_b_10')
// (3, 6, 'neigh_op_bnr_5')
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g0_6')
// (4, 0, 'span4_horz_r_13')
// (4, 0, 'span4_vert_6')
// (4, 1, 'sp4_r_v_b_7')
// (4, 1, 'sp4_v_b_6')
// (4, 1, 'sp4_v_t_47')
// (4, 2, 'sp4_r_v_b_46')
// (4, 2, 'sp4_v_b_47')
// (4, 3, 'sp4_r_v_b_35')
// (4, 3, 'sp4_v_b_34')
// (4, 4, 'neigh_op_top_5')
// (4, 4, 'sp4_r_v_b_22')
// (4, 4, 'sp4_r_v_b_38')
// (4, 4, 'sp4_v_b_23')
// (4, 5, 'lutff_5/out')
// (4, 5, 'sp12_h_r_18')
// (4, 5, 'sp4_r_v_b_11')
// (4, 5, 'sp4_r_v_b_27')
// (4, 5, 'sp4_v_b_10')
// (4, 6, 'neigh_op_bot_5')
// (4, 6, 'sp4_r_v_b_14')
// (4, 7, 'sp4_r_v_b_3')
// (5, 0, 'span4_horz_l_13')
// (5, 0, 'span4_horz_r_1')
// (5, 0, 'span4_vert_7')
// (5, 1, 'sp4_h_r_4')
// (5, 1, 'sp4_v_b_7')
// (5, 1, 'sp4_v_t_46')
// (5, 2, 'sp4_v_b_46')
// (5, 3, 'sp4_h_r_3')
// (5, 3, 'sp4_v_b_35')
// (5, 3, 'sp4_v_t_38')
// (5, 4, 'neigh_op_tnl_5')
// (5, 4, 'sp4_v_b_22')
// (5, 4, 'sp4_v_b_38')
// (5, 5, 'neigh_op_lft_5')
// (5, 5, 'sp12_h_r_21')
// (5, 5, 'sp4_v_b_11')
// (5, 5, 'sp4_v_b_27')
// (5, 6, 'neigh_op_bnl_5')
// (5, 6, 'sp4_v_b_14')
// (5, 7, 'sp4_v_b_3')
// (6, 0, 'io_0/D_OUT_0')
// (6, 0, 'io_0/PAD')
// (6, 0, 'io_1/D_OUT_0')
// (6, 0, 'io_1/PAD')
// (6, 0, 'local_g0_5')
// (6, 0, 'local_g1_5')
// (6, 0, 'span4_horz_r_5')
// (6, 1, 'sp4_h_r_17')
// (6, 3, 'sp4_h_r_14')
// (6, 5, 'sp12_h_r_22')
// (7, 0, 'io_1/D_OUT_0')
// (7, 0, 'io_1/PAD')
// (7, 0, 'local_g0_1')
// (7, 0, 'span12_vert_9')
// (7, 0, 'span4_horz_r_9')
// (7, 1, 'sp12_v_b_9')
// (7, 1, 'sp4_h_r_28')
// (7, 2, 'sp12_v_b_6')
// (7, 3, 'sp12_v_b_5')
// (7, 3, 'sp4_h_r_27')
// (7, 4, 'sp12_v_b_2')
// (7, 5, 'sp12_h_l_22')
// (7, 5, 'sp12_v_b_1')
// (8, 0, 'span4_horz_r_13')
// (8, 1, 'sp4_h_r_41')
// (8, 1, 'sp4_r_v_b_4')
// (8, 3, 'sp4_h_r_38')
// (9, 0, 'io_1/D_OUT_0')
// (9, 0, 'io_1/PAD')
// (9, 0, 'local_g1_4')
// (9, 0, 'span4_horz_l_13')
// (9, 0, 'span4_vert_4')
// (9, 1, 'sp4_h_l_41')
// (9, 1, 'sp4_v_b_4')
// (9, 3, 'sp4_h_l_38')
// (9, 3, 'sp4_h_r_6')
// (10, 0, 'io_0/D_OUT_0')
// (10, 0, 'io_0/PAD')
// (10, 0, 'io_1/D_OUT_0')
// (10, 0, 'io_1/PAD')
// (10, 0, 'local_g0_3')
// (10, 0, 'local_g1_3')
// (10, 0, 'span4_horz_r_3')
// (10, 3, 'sp4_h_r_19')
// (11, 0, 'span4_horz_r_7')
// (11, 3, 'sp4_h_r_30')
// (12, 0, 'span4_horz_r_11')
// (12, 3, 'sp4_h_r_43')
// (13, 1, 'span4_vert_b_11')
// (13, 2, 'span4_vert_b_7')
// (13, 3, 'span4_horz_43')
// (13, 3, 'span4_vert_b_3')

reg n21 = 0;
// (0, 5, 'span4_horz_31')
// (1, 2, 'sp4_r_v_b_42')
// (1, 3, 'neigh_op_tnr_1')
// (1, 3, 'sp4_r_v_b_31')
// (1, 4, 'neigh_op_rgt_1')
// (1, 4, 'sp4_r_v_b_18')
// (1, 5, 'local_g3_2')
// (1, 5, 'lutff_4/in_3')
// (1, 5, 'neigh_op_bnr_1')
// (1, 5, 'sp4_h_r_42')
// (1, 5, 'sp4_r_v_b_7')
// (2, 1, 'sp4_v_t_42')
// (2, 2, 'sp4_v_b_42')
// (2, 3, 'neigh_op_top_1')
// (2, 3, 'sp4_v_b_31')
// (2, 4, 'local_g0_1')
// (2, 4, 'lutff_1/in_2')
// (2, 4, 'lutff_1/out')
// (2, 4, 'sp4_v_b_18')
// (2, 5, 'local_g1_1')
// (2, 5, 'lutff_0/in_0')
// (2, 5, 'lutff_7/in_1')
// (2, 5, 'neigh_op_bot_1')
// (2, 5, 'sp4_h_l_42')
// (2, 5, 'sp4_v_b_7')
// (3, 3, 'neigh_op_tnl_1')
// (3, 4, 'neigh_op_lft_1')
// (3, 5, 'neigh_op_bnl_1')

wire n22;
// (1, 1, 'lutff_7/cout')
// (1, 2, 'carry_in')
// (1, 2, 'carry_in_mux')

reg io_2_0_1 = 0;
// (1, 1, 'sp4_r_v_b_44')
// (1, 2, 'sp4_r_v_b_33')
// (1, 3, 'sp4_r_v_b_20')
// (1, 4, 'sp4_r_v_b_9')
// (2, 0, 'io_1/D_OUT_0')
// (2, 0, 'io_1/PAD')
// (2, 0, 'local_g1_4')
// (2, 0, 'span4_vert_44')
// (2, 1, 'sp4_v_b_44')
// (2, 2, 'sp4_v_b_33')
// (2, 3, 'sp4_v_b_20')
// (2, 4, 'sp4_h_r_9')
// (2, 4, 'sp4_v_b_9')
// (3, 4, 'sp4_h_r_20')
// (4, 4, 'sp4_h_r_33')
// (5, 4, 'sp4_h_r_44')
// (6, 3, 'neigh_op_tnr_2')
// (6, 4, 'neigh_op_rgt_2')
// (6, 4, 'sp4_h_l_44')
// (6, 4, 'sp4_h_r_9')
// (6, 5, 'neigh_op_bnr_2')
// (7, 3, 'neigh_op_top_2')
// (7, 4, 'lutff_2/out')
// (7, 4, 'sp4_h_r_20')
// (7, 5, 'neigh_op_bot_2')
// (8, 3, 'neigh_op_tnl_2')
// (8, 4, 'neigh_op_lft_2')
// (8, 4, 'sp4_h_r_33')
// (8, 5, 'neigh_op_bnl_2')
// (9, 4, 'sp4_h_r_44')
// (10, 4, 'sp4_h_l_44')

wire n24;
// (1, 2, 'local_g2_5')
// (1, 2, 'lutff_4/in_1')
// (1, 2, 'sp4_r_v_b_37')
// (1, 3, 'sp4_r_v_b_24')
// (1, 4, 'neigh_op_tnr_0')
// (1, 4, 'sp4_r_v_b_13')
// (1, 5, 'neigh_op_rgt_0')
// (1, 5, 'sp4_r_v_b_0')
// (1, 6, 'neigh_op_bnr_0')
// (2, 1, 'sp4_v_t_37')
// (2, 2, 'sp4_v_b_37')
// (2, 3, 'sp4_v_b_24')
// (2, 4, 'neigh_op_top_0')
// (2, 4, 'sp4_v_b_13')
// (2, 5, 'lutff_0/out')
// (2, 5, 'sp4_h_r_0')
// (2, 5, 'sp4_v_b_0')
// (2, 6, 'neigh_op_bot_0')
// (3, 4, 'neigh_op_tnl_0')
// (3, 5, 'neigh_op_lft_0')
// (3, 5, 'sp4_h_r_13')
// (3, 6, 'neigh_op_bnl_0')
// (4, 5, 'local_g3_0')
// (4, 5, 'lutff_5/in_0')
// (4, 5, 'sp4_h_r_24')
// (5, 5, 'sp4_h_r_37')
// (6, 5, 'sp4_h_l_37')

reg n25 = 0;
// (1, 2, 'local_g2_6')
// (1, 2, 'lutff_4/in_2')
// (1, 2, 'neigh_op_tnr_6')
// (1, 2, 'sp4_r_v_b_41')
// (1, 3, 'local_g3_6')
// (1, 3, 'lutff_6/in_3')
// (1, 3, 'neigh_op_rgt_6')
// (1, 3, 'sp4_r_v_b_28')
// (1, 4, 'neigh_op_bnr_6')
// (1, 4, 'sp4_r_v_b_17')
// (1, 5, 'sp4_r_v_b_4')
// (2, 1, 'sp4_v_t_41')
// (2, 2, 'neigh_op_top_6')
// (2, 2, 'sp4_r_v_b_40')
// (2, 2, 'sp4_v_b_41')
// (2, 3, 'local_g3_6')
// (2, 3, 'lutff_6/in_1')
// (2, 3, 'lutff_6/out')
// (2, 3, 'sp4_r_v_b_29')
// (2, 3, 'sp4_v_b_28')
// (2, 4, 'neigh_op_bot_6')
// (2, 4, 'sp4_r_v_b_16')
// (2, 4, 'sp4_v_b_17')
// (2, 5, 'local_g0_4')
// (2, 5, 'lutff_7/in_3')
// (2, 5, 'sp4_r_v_b_5')
// (2, 5, 'sp4_v_b_4')
// (3, 1, 'sp4_v_t_40')
// (3, 2, 'neigh_op_tnl_6')
// (3, 2, 'sp4_v_b_40')
// (3, 3, 'neigh_op_lft_6')
// (3, 3, 'sp4_v_b_29')
// (3, 4, 'neigh_op_bnl_6')
// (3, 4, 'sp4_v_b_16')
// (3, 5, 'sp4_h_r_11')
// (3, 5, 'sp4_v_b_5')
// (4, 5, 'local_g0_6')
// (4, 5, 'lutff_5/in_3')
// (4, 5, 'sp4_h_r_22')
// (5, 5, 'sp4_h_r_35')
// (6, 5, 'sp4_h_r_46')
// (7, 5, 'sp4_h_l_46')

reg n26 = 0;
// (1, 2, 'local_g3_7')
// (1, 2, 'lutff_4/in_0')
// (1, 2, 'neigh_op_tnr_7')
// (1, 3, 'local_g3_7')
// (1, 3, 'lutff_7/in_3')
// (1, 3, 'neigh_op_rgt_7')
// (1, 3, 'sp4_r_v_b_46')
// (1, 4, 'neigh_op_bnr_7')
// (1, 4, 'sp4_r_v_b_35')
// (1, 5, 'sp4_r_v_b_22')
// (1, 6, 'sp4_r_v_b_11')
// (2, 2, 'neigh_op_top_7')
// (2, 2, 'sp4_r_v_b_42')
// (2, 2, 'sp4_v_t_46')
// (2, 3, 'local_g0_7')
// (2, 3, 'lutff_7/in_2')
// (2, 3, 'lutff_7/out')
// (2, 3, 'sp4_r_v_b_31')
// (2, 3, 'sp4_v_b_46')
// (2, 4, 'neigh_op_bot_7')
// (2, 4, 'sp4_r_v_b_18')
// (2, 4, 'sp4_v_b_35')
// (2, 5, 'local_g1_6')
// (2, 5, 'lutff_7/in_0')
// (2, 5, 'sp4_r_v_b_7')
// (2, 5, 'sp4_v_b_22')
// (2, 6, 'sp4_v_b_11')
// (3, 1, 'sp4_v_t_42')
// (3, 2, 'neigh_op_tnl_7')
// (3, 2, 'sp4_v_b_42')
// (3, 3, 'neigh_op_lft_7')
// (3, 3, 'sp4_v_b_31')
// (3, 4, 'neigh_op_bnl_7')
// (3, 4, 'sp4_v_b_18')
// (3, 5, 'sp4_h_r_1')
// (3, 5, 'sp4_v_b_7')
// (4, 5, 'local_g0_4')
// (4, 5, 'lutff_5/in_1')
// (4, 5, 'sp4_h_r_12')
// (5, 5, 'sp4_h_r_25')
// (6, 5, 'sp4_h_r_36')
// (7, 5, 'sp4_h_l_36')

wire n27;
// (1, 2, 'lutff_3/cout')
// (1, 2, 'lutff_4/in_3')

reg n28 = 0;
// (1, 2, 'neigh_op_tnr_2')
// (1, 3, 'local_g3_2')
// (1, 3, 'lutff_2/in_3')
// (1, 3, 'neigh_op_rgt_2')
// (1, 4, 'local_g1_2')
// (1, 4, 'lutff_7/in_0')
// (1, 4, 'neigh_op_bnr_2')
// (2, 2, 'neigh_op_top_2')
// (2, 3, 'local_g0_2')
// (2, 3, 'lutff_2/in_2')
// (2, 3, 'lutff_2/out')
// (2, 4, 'local_g1_2')
// (2, 4, 'lutff_5/in_0')
// (2, 4, 'neigh_op_bot_2')
// (3, 2, 'neigh_op_tnl_2')
// (3, 3, 'neigh_op_lft_2')
// (3, 4, 'neigh_op_bnl_2')

reg n29 = 0;
// (1, 2, 'neigh_op_tnr_3')
// (1, 3, 'local_g3_3')
// (1, 3, 'lutff_3/in_3')
// (1, 3, 'neigh_op_rgt_3')
// (1, 4, 'neigh_op_bnr_3')
// (2, 2, 'neigh_op_top_3')
// (2, 3, 'local_g0_3')
// (2, 3, 'lutff_3/in_2')
// (2, 3, 'lutff_3/out')
// (2, 4, 'local_g1_3')
// (2, 4, 'lutff_5/in_1')
// (2, 4, 'lutff_6/in_0')
// (2, 4, 'neigh_op_bot_3')
// (3, 2, 'neigh_op_tnl_3')
// (3, 3, 'neigh_op_lft_3')
// (3, 4, 'neigh_op_bnl_3')

reg n30 = 0;
// (1, 2, 'neigh_op_tnr_4')
// (1, 3, 'local_g3_4')
// (1, 3, 'lutff_4/in_3')
// (1, 3, 'neigh_op_rgt_4')
// (1, 4, 'neigh_op_bnr_4')
// (2, 2, 'neigh_op_top_4')
// (2, 3, 'local_g2_4')
// (2, 3, 'lutff_4/in_2')
// (2, 3, 'lutff_4/out')
// (2, 4, 'local_g0_4')
// (2, 4, 'local_g1_4')
// (2, 4, 'lutff_5/in_3')
// (2, 4, 'lutff_6/in_3')
// (2, 4, 'neigh_op_bot_4')
// (3, 2, 'neigh_op_tnl_4')
// (3, 3, 'neigh_op_lft_4')
// (3, 4, 'neigh_op_bnl_4')

reg n31 = 0;
// (1, 2, 'neigh_op_tnr_5')
// (1, 3, 'local_g3_5')
// (1, 3, 'lutff_5/in_3')
// (1, 3, 'neigh_op_rgt_5')
// (1, 4, 'neigh_op_bnr_5')
// (2, 2, 'neigh_op_top_5')
// (2, 3, 'local_g1_5')
// (2, 3, 'lutff_5/in_1')
// (2, 3, 'lutff_5/out')
// (2, 4, 'local_g0_5')
// (2, 4, 'lutff_6/in_1')
// (2, 4, 'lutff_7/in_2')
// (2, 4, 'neigh_op_bot_5')
// (3, 2, 'neigh_op_tnl_5')
// (3, 3, 'neigh_op_lft_5')
// (3, 4, 'neigh_op_bnl_5')

reg n32 = 0;
// (1, 3, 'local_g2_4')
// (1, 3, 'lutff_1/in_3')
// (1, 3, 'neigh_op_tnr_4')
// (1, 4, 'local_g2_4')
// (1, 4, 'lutff_7/in_1')
// (1, 4, 'neigh_op_rgt_4')
// (1, 5, 'neigh_op_bnr_4')
// (2, 3, 'local_g0_4')
// (2, 3, 'lutff_1/in_1')
// (2, 3, 'neigh_op_top_4')
// (2, 4, 'local_g3_4')
// (2, 4, 'lutff_4/in_3')
// (2, 4, 'lutff_4/out')
// (2, 4, 'lutff_5/in_2')
// (2, 5, 'neigh_op_bot_4')
// (3, 3, 'neigh_op_tnl_4')
// (3, 4, 'neigh_op_lft_4')
// (3, 5, 'neigh_op_bnl_4')

wire n33;
// (1, 3, 'lutff_7/cout')
// (1, 4, 'carry_in')
// (1, 4, 'carry_in_mux')

reg n34 = 0;
// (1, 3, 'neigh_op_tnr_0')
// (1, 4, 'local_g3_0')
// (1, 4, 'lutff_0/in_3')
// (1, 4, 'lutff_7/in_2')
// (1, 4, 'neigh_op_rgt_0')
// (1, 5, 'neigh_op_bnr_0')
// (2, 3, 'neigh_op_top_0')
// (2, 4, 'local_g3_0')
// (2, 4, 'lutff_0/in_1')
// (2, 4, 'lutff_0/out')
// (2, 4, 'lutff_7/in_0')
// (2, 5, 'neigh_op_bot_0')
// (3, 3, 'neigh_op_tnl_0')
// (3, 4, 'neigh_op_lft_0')
// (3, 5, 'neigh_op_bnl_0')

reg n35 = 0;
// (1, 3, 'neigh_op_tnr_2')
// (1, 4, 'local_g3_2')
// (1, 4, 'lutff_2/in_3')
// (1, 4, 'neigh_op_rgt_2')
// (1, 5, 'neigh_op_bnr_2')
// (2, 3, 'neigh_op_top_2')
// (2, 4, 'local_g0_2')
// (2, 4, 'lutff_2/in_2')
// (2, 4, 'lutff_2/out')
// (2, 5, 'local_g1_2')
// (2, 5, 'lutff_0/in_3')
// (2, 5, 'lutff_7/in_2')
// (2, 5, 'neigh_op_bot_2')
// (3, 3, 'neigh_op_tnl_2')
// (3, 4, 'neigh_op_lft_2')
// (3, 5, 'neigh_op_bnl_2')

reg n36 = 0;
// (1, 3, 'neigh_op_tnr_3')
// (1, 4, 'local_g3_3')
// (1, 4, 'lutff_3/in_3')
// (1, 4, 'neigh_op_rgt_3')
// (1, 5, 'neigh_op_bnr_3')
// (2, 3, 'neigh_op_top_3')
// (2, 4, 'local_g3_3')
// (2, 4, 'lutff_3/in_1')
// (2, 4, 'lutff_3/out')
// (2, 4, 'lutff_6/in_2')
// (2, 4, 'lutff_7/in_1')
// (2, 5, 'neigh_op_bot_3')
// (3, 3, 'neigh_op_tnl_3')
// (3, 4, 'neigh_op_lft_3')
// (3, 5, 'neigh_op_bnl_3')

wire n37;
// (1, 3, 'neigh_op_tnr_5')
// (1, 4, 'neigh_op_rgt_5')
// (1, 5, 'neigh_op_bnr_5')
// (2, 3, 'neigh_op_top_5')
// (2, 4, 'lutff_5/out')
// (2, 5, 'local_g1_5')
// (2, 5, 'lutff_0/in_2')
// (2, 5, 'neigh_op_bot_5')
// (3, 3, 'neigh_op_tnl_5')
// (3, 4, 'neigh_op_lft_5')
// (3, 5, 'neigh_op_bnl_5')

wire n38;
// (1, 3, 'neigh_op_tnr_6')
// (1, 4, 'neigh_op_rgt_6')
// (1, 5, 'local_g1_6')
// (1, 5, 'lutff_7/in_0')
// (1, 5, 'neigh_op_bnr_6')
// (2, 3, 'neigh_op_top_6')
// (2, 4, 'lutff_6/out')
// (2, 5, 'neigh_op_bot_6')
// (3, 3, 'neigh_op_tnl_6')
// (3, 4, 'neigh_op_lft_6')
// (3, 5, 'neigh_op_bnl_6')

wire n39;
// (1, 3, 'neigh_op_tnr_7')
// (1, 4, 'neigh_op_rgt_7')
// (1, 5, 'neigh_op_bnr_7')
// (2, 3, 'neigh_op_top_7')
// (2, 4, 'lutff_7/out')
// (2, 5, 'local_g0_7')
// (2, 5, 'lutff_0/in_1')
// (2, 5, 'neigh_op_bot_7')
// (3, 3, 'neigh_op_tnl_7')
// (3, 4, 'neigh_op_lft_7')
// (3, 5, 'neigh_op_bnl_7')

wire n40;
// (1, 4, 'lutff_3/cout')
// (1, 4, 'lutff_4/in_3')

wire n41;
// (1, 4, 'neigh_op_tnr_5')
// (1, 5, 'neigh_op_rgt_5')
// (1, 6, 'neigh_op_bnr_5')
// (2, 4, 'local_g1_5')
// (2, 4, 'lutff_global/s_r')
// (2, 4, 'neigh_op_top_5')
// (2, 5, 'lutff_5/out')
// (2, 6, 'neigh_op_bot_5')
// (3, 4, 'neigh_op_tnl_5')
// (3, 5, 'neigh_op_lft_5')
// (3, 6, 'neigh_op_bnl_5')

wire n42;
// (1, 4, 'neigh_op_tnr_7')
// (1, 5, 'local_g2_7')
// (1, 5, 'lutff_7/in_2')
// (1, 5, 'neigh_op_rgt_7')
// (1, 6, 'neigh_op_bnr_7')
// (2, 4, 'neigh_op_top_7')
// (2, 5, 'lutff_7/out')
// (2, 6, 'neigh_op_bot_7')
// (3, 4, 'neigh_op_tnl_7')
// (3, 5, 'neigh_op_lft_7')
// (3, 6, 'neigh_op_bnl_7')

wire n43;
// (1, 5, 'lutff_6/cout')
// (1, 5, 'lutff_7/in_3')

wire n44;
// (2, 3, 'lutff_1/cout')
// (2, 3, 'lutff_2/in_3')

wire n45;
// (2, 3, 'lutff_2/cout')
// (2, 3, 'lutff_3/in_3')

wire n46;
// (2, 3, 'lutff_3/cout')
// (2, 3, 'lutff_4/in_3')

wire n47;
// (2, 3, 'lutff_4/cout')
// (2, 3, 'lutff_5/in_3')

wire n48;
// (2, 3, 'lutff_5/cout')
// (2, 3, 'lutff_6/in_3')

wire n49;
// (2, 3, 'lutff_6/cout')
// (2, 3, 'lutff_7/in_3')

wire n50;
// (2, 3, 'lutff_7/cout')
// (2, 4, 'carry_in')
// (2, 4, 'carry_in_mux')
// (2, 4, 'lutff_0/in_3')

reg n51 = 0;
// (2, 3, 'sp4_h_r_0')
// (3, 2, 'neigh_op_tnr_4')
// (3, 3, 'neigh_op_rgt_4')
// (3, 3, 'sp4_h_r_13')
// (3, 4, 'neigh_op_bnr_4')
// (4, 2, 'neigh_op_top_4')
// (4, 3, 'local_g1_4')
// (4, 3, 'lutff_4/in_1')
// (4, 3, 'lutff_4/out')
// (4, 3, 'sp4_h_r_24')
// (4, 3, 'sp4_h_r_8')
// (4, 4, 'neigh_op_bot_4')
// (5, 2, 'neigh_op_tnl_4')
// (5, 3, 'neigh_op_lft_4')
// (5, 3, 'sp4_h_r_21')
// (5, 3, 'sp4_h_r_37')
// (5, 4, 'local_g2_4')
// (5, 4, 'lutff_6/in_2')
// (5, 4, 'neigh_op_bnl_4')
// (5, 4, 'sp4_r_v_b_37')
// (5, 5, 'sp4_r_v_b_24')
// (5, 6, 'sp4_r_v_b_13')
// (5, 7, 'sp4_r_v_b_0')
// (6, 3, 'local_g3_0')
// (6, 3, 'lutff_4/in_3')
// (6, 3, 'sp4_h_l_37')
// (6, 3, 'sp4_h_r_32')
// (6, 3, 'sp4_v_t_37')
// (6, 4, 'local_g2_5')
// (6, 4, 'lutff_7/in_0')
// (6, 4, 'sp4_v_b_37')
// (6, 5, 'sp4_v_b_24')
// (6, 6, 'sp4_v_b_13')
// (6, 7, 'sp4_v_b_0')
// (7, 3, 'sp4_h_r_45')
// (8, 3, 'sp4_h_l_45')

reg n52 = 0;
// (2, 3, 'sp4_h_r_2')
// (3, 2, 'neigh_op_tnr_5')
// (3, 3, 'neigh_op_rgt_5')
// (3, 3, 'sp4_h_r_15')
// (3, 4, 'neigh_op_bnr_5')
// (4, 2, 'neigh_op_top_5')
// (4, 3, 'local_g3_5')
// (4, 3, 'lutff_5/in_1')
// (4, 3, 'lutff_5/out')
// (4, 3, 'sp4_h_r_10')
// (4, 3, 'sp4_h_r_26')
// (4, 4, 'neigh_op_bot_5')
// (5, 2, 'neigh_op_tnl_5')
// (5, 3, 'neigh_op_lft_5')
// (5, 3, 'sp4_h_r_23')
// (5, 3, 'sp4_h_r_39')
// (5, 4, 'local_g3_5')
// (5, 4, 'lutff_7/in_1')
// (5, 4, 'neigh_op_bnl_5')
// (5, 4, 'sp4_r_v_b_42')
// (5, 5, 'sp4_r_v_b_31')
// (5, 6, 'sp4_r_v_b_18')
// (5, 7, 'sp4_r_v_b_7')
// (6, 3, 'sp4_h_l_39')
// (6, 3, 'sp4_h_r_34')
// (6, 3, 'sp4_v_t_42')
// (6, 4, 'local_g3_2')
// (6, 4, 'lutff_7/in_2')
// (6, 4, 'sp4_v_b_42')
// (6, 5, 'sp4_v_b_31')
// (6, 6, 'sp4_v_b_18')
// (6, 7, 'sp4_v_b_7')
// (7, 3, 'local_g3_7')
// (7, 3, 'lutff_3/in_3')
// (7, 3, 'sp4_h_r_47')
// (8, 3, 'sp4_h_l_47')

wire n53;
// (2, 4, 'lutff_0/cout')
// (2, 4, 'lutff_1/in_3')

wire n54;
// (2, 4, 'lutff_1/cout')
// (2, 4, 'lutff_2/in_3')

wire n55;
// (2, 4, 'lutff_2/cout')
// (2, 4, 'lutff_3/in_3')

reg n56 = 0;
// (3, 2, 'neigh_op_tnr_2')
// (3, 3, 'neigh_op_rgt_2')
// (3, 4, 'neigh_op_bnr_2')
// (4, 2, 'neigh_op_top_2')
// (4, 3, 'local_g2_2')
// (4, 3, 'lutff_2/in_2')
// (4, 3, 'lutff_2/out')
// (4, 4, 'local_g1_2')
// (4, 4, 'lutff_5/in_0')
// (4, 4, 'neigh_op_bot_2')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'local_g1_2')
// (5, 3, 'lutff_2/in_3')
// (5, 3, 'neigh_op_lft_2')
// (5, 4, 'local_g3_2')
// (5, 4, 'lutff_5/in_2')
// (5, 4, 'lutff_7/in_0')
// (5, 4, 'neigh_op_bnl_2')

reg n57 = 0;
// (3, 2, 'neigh_op_tnr_3')
// (3, 3, 'neigh_op_rgt_3')
// (3, 4, 'neigh_op_bnr_3')
// (4, 2, 'neigh_op_top_3')
// (4, 3, 'local_g1_3')
// (4, 3, 'lutff_3/in_1')
// (4, 3, 'lutff_3/out')
// (4, 4, 'local_g1_3')
// (4, 4, 'lutff_5/in_1')
// (4, 4, 'neigh_op_bot_3')
// (5, 2, 'neigh_op_tnl_3')
// (5, 3, 'local_g1_3')
// (5, 3, 'lutff_3/in_3')
// (5, 3, 'neigh_op_lft_3')
// (5, 4, 'local_g2_3')
// (5, 4, 'local_g3_3')
// (5, 4, 'lutff_5/in_1')
// (5, 4, 'lutff_7/in_2')
// (5, 4, 'neigh_op_bnl_3')

reg n58 = 0;
// (3, 2, 'neigh_op_tnr_6')
// (3, 3, 'neigh_op_rgt_6')
// (3, 3, 'sp4_h_r_1')
// (3, 4, 'neigh_op_bnr_6')
// (4, 1, 'sp4_r_v_b_37')
// (4, 2, 'neigh_op_top_6')
// (4, 2, 'sp4_r_v_b_24')
// (4, 3, 'local_g1_6')
// (4, 3, 'lutff_6/in_1')
// (4, 3, 'lutff_6/out')
// (4, 3, 'sp4_h_r_12')
// (4, 3, 'sp4_r_v_b_13')
// (4, 4, 'neigh_op_bot_6')
// (4, 4, 'sp4_r_v_b_0')
// (5, 0, 'span4_vert_37')
// (5, 1, 'sp4_v_b_37')
// (5, 2, 'neigh_op_tnl_6')
// (5, 2, 'sp4_v_b_24')
// (5, 3, 'neigh_op_lft_6')
// (5, 3, 'sp4_h_r_25')
// (5, 3, 'sp4_v_b_13')
// (5, 4, 'local_g2_6')
// (5, 4, 'lutff_6/in_0')
// (5, 4, 'neigh_op_bnl_6')
// (5, 4, 'sp4_h_r_6')
// (5, 4, 'sp4_v_b_0')
// (6, 3, 'local_g3_4')
// (6, 3, 'lutff_6/in_3')
// (6, 3, 'sp4_h_r_36')
// (6, 4, 'local_g1_3')
// (6, 4, 'lutff_7/in_1')
// (6, 4, 'sp4_h_r_19')
// (7, 3, 'sp4_h_l_36')
// (7, 4, 'sp4_h_r_30')
// (8, 4, 'sp4_h_r_43')
// (9, 4, 'sp4_h_l_43')

reg n59 = 0;
// (3, 2, 'neigh_op_tnr_7')
// (3, 3, 'neigh_op_rgt_7')
// (3, 3, 'sp4_h_r_3')
// (3, 4, 'neigh_op_bnr_7')
// (4, 1, 'sp4_r_v_b_39')
// (4, 2, 'neigh_op_top_7')
// (4, 2, 'sp4_r_v_b_26')
// (4, 3, 'local_g1_7')
// (4, 3, 'lutff_7/in_1')
// (4, 3, 'lutff_7/out')
// (4, 3, 'sp4_h_r_14')
// (4, 3, 'sp4_r_v_b_15')
// (4, 4, 'neigh_op_bot_7')
// (4, 4, 'sp4_r_v_b_2')
// (5, 0, 'span4_vert_39')
// (5, 1, 'sp4_v_b_39')
// (5, 2, 'neigh_op_tnl_7')
// (5, 2, 'sp4_v_b_26')
// (5, 3, 'neigh_op_lft_7')
// (5, 3, 'sp4_h_r_27')
// (5, 3, 'sp4_v_b_15')
// (5, 4, 'local_g2_7')
// (5, 4, 'lutff_6/in_3')
// (5, 4, 'neigh_op_bnl_7')
// (5, 4, 'sp4_h_r_2')
// (5, 4, 'sp4_v_b_2')
// (6, 3, 'local_g2_6')
// (6, 3, 'lutff_7/in_3')
// (6, 3, 'sp4_h_r_38')
// (6, 4, 'local_g1_7')
// (6, 4, 'lutff_7/in_3')
// (6, 4, 'sp4_h_r_15')
// (7, 3, 'sp4_h_l_38')
// (7, 4, 'sp4_h_r_26')
// (8, 4, 'sp4_h_r_39')
// (9, 4, 'sp4_h_l_39')

reg n60 = 0;
// (3, 3, 'neigh_op_tnr_0')
// (3, 4, 'neigh_op_rgt_0')
// (3, 5, 'neigh_op_bnr_0')
// (4, 3, 'neigh_op_top_0')
// (4, 4, 'local_g2_0')
// (4, 4, 'lutff_0/in_2')
// (4, 4, 'lutff_0/out')
// (4, 4, 'lutff_7/in_3')
// (4, 4, 'sp4_h_r_0')
// (4, 5, 'neigh_op_bot_0')
// (5, 3, 'neigh_op_tnl_0')
// (5, 4, 'local_g1_0')
// (5, 4, 'lutff_6/in_1')
// (5, 4, 'neigh_op_lft_0')
// (5, 4, 'sp4_h_r_13')
// (5, 5, 'neigh_op_bnl_0')
// (6, 4, 'local_g3_0')
// (6, 4, 'lutff_0/in_3')
// (6, 4, 'sp4_h_r_24')
// (7, 4, 'sp4_h_r_37')
// (8, 4, 'sp4_h_l_37')

reg n61 = 0;
// (3, 3, 'neigh_op_tnr_1')
// (3, 4, 'neigh_op_rgt_1')
// (3, 5, 'neigh_op_bnr_1')
// (4, 3, 'neigh_op_top_1')
// (4, 4, 'local_g0_1')
// (4, 4, 'lutff_1/in_2')
// (4, 4, 'lutff_1/out')
// (4, 4, 'lutff_7/in_2')
// (4, 4, 'sp4_h_r_2')
// (4, 5, 'neigh_op_bot_1')
// (5, 3, 'neigh_op_tnl_1')
// (5, 4, 'local_g1_1')
// (5, 4, 'lutff_7/in_3')
// (5, 4, 'neigh_op_lft_1')
// (5, 4, 'sp4_h_r_15')
// (5, 5, 'neigh_op_bnl_1')
// (6, 4, 'local_g2_2')
// (6, 4, 'lutff_1/in_3')
// (6, 4, 'sp4_h_r_26')
// (7, 4, 'sp4_h_r_39')
// (8, 4, 'sp4_h_l_39')

reg n62 = 0;
// (3, 3, 'neigh_op_tnr_2')
// (3, 4, 'neigh_op_rgt_2')
// (3, 5, 'neigh_op_bnr_2')
// (4, 3, 'neigh_op_top_2')
// (4, 4, 'local_g0_2')
// (4, 4, 'lutff_2/in_2')
// (4, 4, 'lutff_2/out')
// (4, 4, 'lutff_7/in_1')
// (4, 4, 'sp4_h_r_4')
// (4, 5, 'neigh_op_bot_2')
// (5, 3, 'neigh_op_tnl_2')
// (5, 4, 'neigh_op_lft_2')
// (5, 4, 'sp4_h_r_17')
// (5, 5, 'local_g2_2')
// (5, 5, 'lutff_7/in_1')
// (5, 5, 'neigh_op_bnl_2')
// (6, 4, 'sp4_h_r_28')
// (7, 4, 'local_g2_1')
// (7, 4, 'lutff_0/in_3')
// (7, 4, 'sp4_h_r_41')
// (8, 4, 'sp4_h_l_41')

reg n63 = 0;
// (3, 3, 'neigh_op_tnr_3')
// (3, 4, 'neigh_op_rgt_3')
// (3, 5, 'neigh_op_bnr_3')
// (4, 3, 'neigh_op_top_3')
// (4, 4, 'local_g2_3')
// (4, 4, 'lutff_3/in_0')
// (4, 4, 'lutff_3/out')
// (4, 4, 'lutff_7/in_0')
// (4, 4, 'sp4_h_r_6')
// (4, 5, 'neigh_op_bot_3')
// (5, 3, 'neigh_op_tnl_3')
// (5, 4, 'neigh_op_lft_3')
// (5, 4, 'sp4_h_r_19')
// (5, 5, 'local_g3_3')
// (5, 5, 'lutff_7/in_3')
// (5, 5, 'neigh_op_bnl_3')
// (6, 4, 'sp4_h_r_30')
// (7, 4, 'local_g3_3')
// (7, 4, 'lutff_1/in_3')
// (7, 4, 'sp4_h_r_43')
// (8, 4, 'sp4_h_l_43')

wire n64;
// (3, 3, 'neigh_op_tnr_5')
// (3, 4, 'neigh_op_rgt_5')
// (3, 5, 'neigh_op_bnr_5')
// (4, 3, 'neigh_op_top_5')
// (4, 4, 'lutff_5/out')
// (4, 5, 'neigh_op_bot_5')
// (5, 3, 'neigh_op_tnl_5')
// (5, 4, 'local_g1_5')
// (5, 4, 'lutff_4/in_0')
// (5, 4, 'neigh_op_lft_5')
// (5, 5, 'neigh_op_bnl_5')

reg n65 = 0;
// (3, 3, 'neigh_op_tnr_6')
// (3, 4, 'neigh_op_rgt_6')
// (3, 5, 'neigh_op_bnr_6')
// (4, 3, 'local_g0_6')
// (4, 3, 'lutff_1/in_1')
// (4, 3, 'neigh_op_top_6')
// (4, 4, 'local_g0_6')
// (4, 4, 'lutff_5/in_3')
// (4, 4, 'lutff_6/in_2')
// (4, 4, 'lutff_6/out')
// (4, 5, 'neigh_op_bot_6')
// (5, 3, 'local_g2_6')
// (5, 3, 'lutff_1/in_3')
// (5, 3, 'neigh_op_tnl_6')
// (5, 4, 'local_g1_6')
// (5, 4, 'lutff_5/in_0')
// (5, 4, 'neigh_op_lft_6')
// (5, 5, 'local_g3_6')
// (5, 5, 'lutff_7/in_0')
// (5, 5, 'neigh_op_bnl_6')

wire n66;
// (3, 3, 'neigh_op_tnr_7')
// (3, 4, 'neigh_op_rgt_7')
// (3, 4, 'sp4_h_r_3')
// (3, 5, 'neigh_op_bnr_7')
// (4, 3, 'neigh_op_top_7')
// (4, 4, 'lutff_7/out')
// (4, 4, 'sp4_h_r_14')
// (4, 5, 'neigh_op_bot_7')
// (5, 3, 'neigh_op_tnl_7')
// (5, 4, 'local_g0_7')
// (5, 4, 'lutff_4/in_1')
// (5, 4, 'neigh_op_lft_7')
// (5, 4, 'sp4_h_r_27')
// (5, 5, 'neigh_op_bnl_7')
// (6, 4, 'sp4_h_r_38')
// (7, 4, 'local_g0_6')
// (7, 4, 'lutff_2/in_2')
// (7, 4, 'sp4_h_l_38')
// (7, 4, 'sp4_h_r_6')
// (8, 4, 'sp4_h_r_19')
// (9, 4, 'sp4_h_r_30')
// (10, 4, 'sp4_h_r_43')
// (11, 4, 'sp4_h_l_43')

wire n67;
// (3, 4, 'sp4_h_r_2')
// (4, 3, 'neigh_op_tnr_5')
// (4, 4, 'neigh_op_rgt_5')
// (4, 4, 'sp4_h_r_15')
// (4, 5, 'neigh_op_bnr_5')
// (5, 3, 'neigh_op_top_5')
// (5, 4, 'lutff_5/out')
// (5, 4, 'sp4_h_r_26')
// (5, 5, 'neigh_op_bot_5')
// (6, 3, 'neigh_op_tnl_5')
// (6, 4, 'neigh_op_lft_5')
// (6, 4, 'sp4_h_r_39')
// (6, 5, 'neigh_op_bnl_5')
// (7, 4, 'local_g0_2')
// (7, 4, 'lutff_2/in_0')
// (7, 4, 'sp4_h_l_39')
// (7, 4, 'sp4_h_r_2')
// (8, 4, 'sp4_h_r_15')
// (9, 4, 'sp4_h_r_26')
// (10, 4, 'sp4_h_r_39')
// (11, 4, 'sp4_h_l_39')

wire n68;
// (4, 2, 'neigh_op_tnr_1')
// (4, 3, 'neigh_op_rgt_1')
// (4, 4, 'neigh_op_bnr_1')
// (5, 2, 'neigh_op_top_1')
// (5, 3, 'local_g2_1')
// (5, 3, 'lutff_1/in_2')
// (5, 3, 'lutff_1/out')
// (5, 4, 'neigh_op_bot_1')
// (6, 2, 'neigh_op_tnl_1')
// (6, 3, 'local_g1_1')
// (6, 3, 'lutff_1/in_1')
// (6, 3, 'neigh_op_lft_1')
// (6, 4, 'neigh_op_bnl_1')

wire n69;
// (4, 2, 'neigh_op_tnr_2')
// (4, 3, 'neigh_op_rgt_2')
// (4, 4, 'neigh_op_bnr_2')
// (5, 2, 'neigh_op_top_2')
// (5, 3, 'local_g0_2')
// (5, 3, 'lutff_2/in_2')
// (5, 3, 'lutff_2/out')
// (5, 3, 'sp4_h_r_4')
// (5, 4, 'neigh_op_bot_2')
// (6, 2, 'neigh_op_tnl_2')
// (6, 3, 'local_g1_2')
// (6, 3, 'lutff_2/in_1')
// (6, 3, 'neigh_op_lft_2')
// (6, 3, 'sp4_h_r_17')
// (6, 4, 'neigh_op_bnl_2')
// (7, 3, 'local_g3_4')
// (7, 3, 'lutff_0/in_1')
// (7, 3, 'sp4_h_r_28')
// (8, 3, 'sp4_h_r_41')
// (9, 3, 'sp4_h_l_41')

wire n70;
// (4, 2, 'neigh_op_tnr_3')
// (4, 3, 'neigh_op_rgt_3')
// (4, 4, 'neigh_op_bnr_3')
// (5, 2, 'neigh_op_top_3')
// (5, 3, 'local_g2_3')
// (5, 3, 'lutff_3/in_2')
// (5, 3, 'lutff_3/out')
// (5, 3, 'sp4_h_r_6')
// (5, 4, 'neigh_op_bot_3')
// (6, 2, 'neigh_op_tnl_3')
// (6, 3, 'local_g1_3')
// (6, 3, 'lutff_3/in_1')
// (6, 3, 'neigh_op_lft_3')
// (6, 3, 'sp4_h_r_19')
// (6, 4, 'neigh_op_bnl_3')
// (7, 3, 'local_g2_6')
// (7, 3, 'lutff_1/in_1')
// (7, 3, 'sp4_h_r_30')
// (8, 3, 'sp4_h_r_43')
// (9, 3, 'sp4_h_l_43')

reg n71 = 0;
// (4, 2, 'sp4_r_v_b_45')
// (4, 3, 'local_g2_0')
// (4, 3, 'lutff_0/in_2')
// (4, 3, 'sp4_r_v_b_32')
// (4, 4, 'local_g3_4')
// (4, 4, 'lutff_5/in_2')
// (4, 4, 'lutff_6/in_3')
// (4, 4, 'neigh_op_tnr_4')
// (4, 4, 'sp4_r_v_b_21')
// (4, 5, 'neigh_op_rgt_4')
// (4, 5, 'sp4_r_v_b_8')
// (4, 6, 'neigh_op_bnr_4')
// (5, 1, 'sp4_v_t_45')
// (5, 2, 'sp4_v_b_45')
// (5, 3, 'sp4_v_b_32')
// (5, 4, 'local_g0_4')
// (5, 4, 'lutff_5/in_3')
// (5, 4, 'neigh_op_top_4')
// (5, 4, 'sp4_v_b_21')
// (5, 5, 'local_g3_4')
// (5, 5, 'lutff_4/out')
// (5, 5, 'lutff_7/in_2')
// (5, 5, 'sp4_v_b_8')
// (5, 6, 'neigh_op_bot_4')
// (6, 4, 'local_g3_4')
// (6, 4, 'lutff_5/in_0')
// (6, 4, 'neigh_op_tnl_4')
// (6, 5, 'neigh_op_lft_4')
// (6, 6, 'neigh_op_bnl_4')

wire n72;
// (4, 3, 'local_g2_4')
// (4, 3, 'lutff_global/s_r')
// (4, 3, 'neigh_op_tnr_4')
// (4, 4, 'local_g2_4')
// (4, 4, 'lutff_global/s_r')
// (4, 4, 'neigh_op_rgt_4')
// (4, 5, 'neigh_op_bnr_4')
// (5, 3, 'neigh_op_top_4')
// (5, 4, 'lutff_4/out')
// (5, 5, 'local_g0_4')
// (5, 5, 'lutff_global/s_r')
// (5, 5, 'neigh_op_bot_4')
// (6, 3, 'neigh_op_tnl_4')
// (6, 4, 'neigh_op_lft_4')
// (6, 5, 'neigh_op_bnl_4')

wire n73;
// (4, 3, 'lutff_1/cout')
// (4, 3, 'lutff_2/in_3')

wire n74;
// (4, 3, 'lutff_2/cout')
// (4, 3, 'lutff_3/in_3')

wire n75;
// (4, 3, 'lutff_3/cout')
// (4, 3, 'lutff_4/in_3')

wire n76;
// (4, 3, 'lutff_4/cout')
// (4, 3, 'lutff_5/in_3')

wire n77;
// (4, 3, 'lutff_5/cout')
// (4, 3, 'lutff_6/in_3')

wire n78;
// (4, 3, 'lutff_6/cout')
// (4, 3, 'lutff_7/in_3')

wire n79;
// (4, 3, 'lutff_7/cout')
// (4, 4, 'carry_in')
// (4, 4, 'carry_in_mux')
// (4, 4, 'lutff_0/in_3')

wire n80;
// (4, 3, 'neigh_op_tnr_6')
// (4, 4, 'neigh_op_rgt_6')
// (4, 5, 'neigh_op_bnr_6')
// (5, 3, 'neigh_op_top_6')
// (5, 4, 'lutff_6/out')
// (5, 5, 'local_g0_6')
// (5, 5, 'lutff_3/in_3')
// (5, 5, 'neigh_op_bot_6')
// (6, 3, 'neigh_op_tnl_6')
// (6, 4, 'neigh_op_lft_6')
// (6, 5, 'neigh_op_bnl_6')

wire n81;
// (4, 3, 'neigh_op_tnr_7')
// (4, 4, 'neigh_op_rgt_7')
// (4, 5, 'neigh_op_bnr_7')
// (5, 3, 'neigh_op_top_7')
// (5, 4, 'lutff_7/out')
// (5, 5, 'local_g0_7')
// (5, 5, 'lutff_3/in_2')
// (5, 5, 'neigh_op_bot_7')
// (6, 3, 'neigh_op_tnl_7')
// (6, 4, 'neigh_op_lft_7')
// (6, 5, 'neigh_op_bnl_7')

wire n82;
// (4, 3, 'sp4_h_r_3')
// (5, 3, 'local_g1_6')
// (5, 3, 'lutff_5/in_2')
// (5, 3, 'sp4_h_r_14')
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'local_g2_3')
// (6, 3, 'lutff_5/in_2')
// (6, 3, 'neigh_op_rgt_3')
// (6, 3, 'sp4_h_r_27')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'local_g2_3')
// (7, 3, 'lutff_3/in_2')
// (7, 3, 'lutff_3/out')
// (7, 3, 'sp4_h_r_38')
// (7, 4, 'neigh_op_bot_3')
// (8, 2, 'neigh_op_tnl_3')
// (8, 3, 'neigh_op_lft_3')
// (8, 3, 'sp4_h_l_38')
// (8, 4, 'neigh_op_bnl_3')

wire n83;
// (4, 4, 'lutff_0/cout')
// (4, 4, 'lutff_1/in_3')

wire n84;
// (4, 4, 'lutff_1/cout')
// (4, 4, 'lutff_2/in_3')

wire n85;
// (4, 4, 'lutff_2/cout')
// (4, 4, 'lutff_3/in_3')

wire n86;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'local_g2_3')
// (4, 5, 'lutff_5/in_2')
// (4, 5, 'neigh_op_rgt_3')
// (4, 6, 'neigh_op_bnr_3')
// (5, 4, 'neigh_op_top_3')
// (5, 5, 'lutff_3/out')
// (5, 6, 'neigh_op_bot_3')
// (6, 4, 'neigh_op_tnl_3')
// (6, 5, 'neigh_op_lft_3')
// (6, 6, 'neigh_op_bnl_3')

wire n87;
// (4, 4, 'neigh_op_tnr_7')
// (4, 5, 'neigh_op_rgt_7')
// (4, 6, 'neigh_op_bnr_7')
// (5, 4, 'neigh_op_top_7')
// (5, 5, 'local_g1_7')
// (5, 5, 'lutff_3/in_1')
// (5, 5, 'lutff_7/out')
// (5, 6, 'neigh_op_bot_7')
// (6, 4, 'neigh_op_tnl_7')
// (6, 5, 'neigh_op_lft_7')
// (6, 6, 'neigh_op_bnl_7')

wire n88;
// (5, 2, 'neigh_op_tnr_4')
// (5, 3, 'local_g2_4')
// (5, 3, 'lutff_4/in_2')
// (5, 3, 'neigh_op_rgt_4')
// (5, 4, 'neigh_op_bnr_4')
// (6, 2, 'neigh_op_top_4')
// (6, 3, 'local_g1_4')
// (6, 3, 'lutff_4/in_1')
// (6, 3, 'lutff_4/out')
// (6, 4, 'neigh_op_bot_4')
// (7, 2, 'neigh_op_tnl_4')
// (7, 3, 'local_g0_4')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'neigh_op_lft_4')
// (7, 4, 'neigh_op_bnl_4')

wire n89;
// (5, 2, 'neigh_op_tnr_6')
// (5, 3, 'local_g3_6')
// (5, 3, 'lutff_6/in_1')
// (5, 3, 'neigh_op_rgt_6')
// (5, 4, 'neigh_op_bnr_6')
// (6, 2, 'neigh_op_top_6')
// (6, 3, 'local_g3_6')
// (6, 3, 'lutff_6/in_1')
// (6, 3, 'lutff_6/out')
// (6, 4, 'neigh_op_bot_6')
// (7, 2, 'neigh_op_tnl_6')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_4/in_1')
// (7, 3, 'neigh_op_lft_6')
// (7, 4, 'neigh_op_bnl_6')

wire n90;
// (5, 2, 'neigh_op_tnr_7')
// (5, 3, 'local_g3_7')
// (5, 3, 'lutff_7/in_1')
// (5, 3, 'neigh_op_rgt_7')
// (5, 4, 'neigh_op_bnr_7')
// (6, 2, 'neigh_op_top_7')
// (6, 3, 'local_g0_7')
// (6, 3, 'lutff_7/in_2')
// (6, 3, 'lutff_7/out')
// (6, 4, 'neigh_op_bot_7')
// (7, 2, 'neigh_op_tnl_7')
// (7, 3, 'local_g1_7')
// (7, 3, 'lutff_5/in_1')
// (7, 3, 'neigh_op_lft_7')
// (7, 4, 'neigh_op_bnl_7')

wire n91;
// (5, 3, 'local_g2_5')
// (5, 3, 'lutff_0/in_1')
// (5, 3, 'neigh_op_tnr_5')
// (5, 4, 'neigh_op_rgt_5')
// (5, 5, 'local_g1_5')
// (5, 5, 'lutff_4/in_0')
// (5, 5, 'neigh_op_bnr_5')
// (6, 3, 'local_g0_5')
// (6, 3, 'lutff_0/in_1')
// (6, 3, 'neigh_op_top_5')
// (6, 4, 'lutff_5/out')
// (6, 5, 'neigh_op_bot_5')
// (7, 3, 'neigh_op_tnl_5')
// (7, 4, 'neigh_op_lft_5')
// (7, 5, 'neigh_op_bnl_5')

wire n92;
// (5, 3, 'lutff_7/cout')
// (5, 4, 'carry_in')
// (5, 4, 'carry_in_mux')

wire n93;
// (5, 3, 'neigh_op_tnr_0')
// (5, 4, 'local_g3_0')
// (5, 4, 'lutff_0/in_1')
// (5, 4, 'neigh_op_rgt_0')
// (5, 5, 'neigh_op_bnr_0')
// (6, 3, 'neigh_op_top_0')
// (6, 4, 'local_g0_0')
// (6, 4, 'lutff_0/in_2')
// (6, 4, 'lutff_0/out')
// (6, 5, 'neigh_op_bot_0')
// (7, 3, 'local_g2_0')
// (7, 3, 'lutff_6/in_2')
// (7, 3, 'neigh_op_tnl_0')
// (7, 4, 'neigh_op_lft_0')
// (7, 5, 'neigh_op_bnl_0')

wire n94;
// (5, 3, 'neigh_op_tnr_1')
// (5, 4, 'local_g2_1')
// (5, 4, 'lutff_1/in_2')
// (5, 4, 'neigh_op_rgt_1')
// (5, 5, 'neigh_op_bnr_1')
// (6, 3, 'neigh_op_top_1')
// (6, 4, 'local_g0_1')
// (6, 4, 'lutff_1/in_2')
// (6, 4, 'lutff_1/out')
// (6, 5, 'neigh_op_bot_1')
// (7, 3, 'local_g3_1')
// (7, 3, 'lutff_7/in_1')
// (7, 3, 'neigh_op_tnl_1')
// (7, 4, 'neigh_op_lft_1')
// (7, 5, 'neigh_op_bnl_1')

wire n95;
// (5, 3, 'neigh_op_tnr_4')
// (5, 4, 'neigh_op_rgt_4')
// (5, 5, 'local_g1_4')
// (5, 5, 'lutff_3/in_0')
// (5, 5, 'neigh_op_bnr_4')
// (6, 3, 'neigh_op_top_4')
// (6, 4, 'lutff_4/out')
// (6, 5, 'neigh_op_bot_4')
// (7, 3, 'neigh_op_tnl_4')
// (7, 4, 'neigh_op_lft_4')
// (7, 5, 'neigh_op_bnl_4')

wire n96;
// (5, 3, 'neigh_op_tnr_7')
// (5, 4, 'local_g3_7')
// (5, 4, 'lutff_4/in_2')
// (5, 4, 'neigh_op_rgt_7')
// (5, 5, 'neigh_op_bnr_7')
// (6, 3, 'neigh_op_top_7')
// (6, 4, 'lutff_7/out')
// (6, 5, 'neigh_op_bot_7')
// (7, 3, 'neigh_op_tnl_7')
// (7, 4, 'local_g0_7')
// (7, 4, 'lutff_2/in_1')
// (7, 4, 'neigh_op_lft_7')
// (7, 5, 'neigh_op_bnl_7')

wire n97;
// (5, 4, 'local_g0_0')
// (5, 4, 'lutff_2/in_2')
// (5, 4, 'sp4_h_r_8')
// (6, 3, 'neigh_op_tnr_0')
// (6, 4, 'local_g2_0')
// (6, 4, 'lutff_2/in_2')
// (6, 4, 'neigh_op_rgt_0')
// (6, 4, 'sp4_h_r_21')
// (6, 5, 'neigh_op_bnr_0')
// (7, 3, 'neigh_op_top_0')
// (7, 4, 'local_g1_0')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'lutff_0/out')
// (7, 4, 'sp4_h_r_32')
// (7, 5, 'neigh_op_bot_0')
// (8, 3, 'neigh_op_tnl_0')
// (8, 4, 'neigh_op_lft_0')
// (8, 4, 'sp4_h_r_45')
// (8, 5, 'neigh_op_bnl_0')
// (9, 4, 'sp4_h_l_45')

wire n98;
// (5, 4, 'local_g1_2')
// (5, 4, 'lutff_3/in_2')
// (5, 4, 'sp4_h_r_10')
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'local_g2_1')
// (6, 4, 'lutff_3/in_2')
// (6, 4, 'neigh_op_rgt_1')
// (6, 4, 'sp4_h_r_23')
// (6, 5, 'neigh_op_bnr_1')
// (7, 3, 'neigh_op_top_1')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_1/in_2')
// (7, 4, 'lutff_1/out')
// (7, 4, 'sp4_h_r_34')
// (7, 5, 'neigh_op_bot_1')
// (8, 3, 'neigh_op_tnl_1')
// (8, 4, 'neigh_op_lft_1')
// (8, 4, 'sp4_h_r_47')
// (8, 5, 'neigh_op_bnl_1')
// (9, 4, 'sp4_h_l_47')

wire n99;
// (5, 4, 'lutff_3/cout')
// (5, 4, 'lutff_4/in_3')

wire n100;
// (6, 3, 'lutff_7/cout')
// (6, 4, 'carry_in')
// (6, 4, 'carry_in_mux')

wire n101;
// (6, 4, 'lutff_3/cout')
// (6, 4, 'lutff_4/in_3')

wire n102;
// (7, 3, 'lutff_7/cout')
// (7, 4, 'carry_in')
// (7, 4, 'carry_in_mux')

wire n103;
// (7, 4, 'lutff_1/cout')
// (7, 4, 'lutff_2/in_3')

wire n104;
// (5, 3, 'lutff_3/cout')

wire n105;
// (5, 4, 'lutff_2/cout')

wire n106;
// (7, 3, 'lutff_5/cout')

wire n107;
// (1, 3, 'lutff_0/cout')

wire n108;
// (1, 1, 'lutff_0/cout')

wire n109;
// (5, 3, 'lutff_5/cout')

wire n110;
// (1, 5, 'lutff_0/cout')

wire n111;
// (1, 3, 'lutff_2/cout')

wire n112;
// (1, 1, 'lutff_2/cout')

wire n113;
// (7, 3, 'lutff_0/cout')

wire n114;
// (1, 5, 'lutff_2/cout')

wire n115;
// (1, 3, 'lutff_4/cout')

wire n116;
// (1, 1, 'lutff_4/cout')

wire n117;
// (5, 3, 'lutff_0/cout')

wire n118;
// (7, 3, 'lutff_2/cout')

wire n119;
// (1, 5, 'lutff_4/cout')

wire n120;
// (1, 3, 'lutff_6/cout')

wire n121;
// (5, 3, 'lutff_2/cout')

wire n122;
// (5, 4, 'lutff_1/cout')

wire n123;
// (7, 3, 'lutff_4/cout')

wire n124;
// (6, 3, 'lutff_1/cout')

wire n125;
// (1, 2, 'lutff_1/cout')

wire n126;
// (6, 3, 'lutff_3/cout')

wire n127;
// (1, 3, 'lutff_1/cout')

wire n128;
// (1, 4, 'lutff_0/cout')

wire n129;
// (6, 4, 'lutff_1/cout')

wire n130;
// (1, 5, 'lutff_1/cout')

wire n131;
// (6, 3, 'lutff_5/cout')

wire n132;
// (1, 3, 'lutff_3/cout')

wire n133;
// (1, 4, 'lutff_2/cout')

wire n134;
// (7, 4, 'lutff_0/cout')

wire n135;
// (1, 1, 'lutff_6/cout')

wire n136;
// (1, 4, 'lutff_4/cout')

wire n137;
// (5, 4, 'lutff_0/cout')

wire n138;
// (5, 3, 'lutff_4/cout')

wire n139;
// (7, 3, 'lutff_6/cout')

wire n140;
// (6, 3, 'lutff_0/cout')

wire n141;
// (1, 2, 'lutff_0/cout')

wire n142;
// (4, 3, 'lutff_0/cout')

wire n143;
// (1, 1, 'lutff_1/cout')

wire n144;
// (5, 3, 'lutff_6/cout')

wire n145;
// (6, 3, 'lutff_2/cout')

wire n146;
// (1, 2, 'lutff_2/cout')

wire n147;
// (2, 3, 'lutff_0/cout')

wire n148;
// (6, 4, 'lutff_0/cout')

wire n149;
// (1, 1, 'lutff_3/cout')

wire n150;
// (7, 3, 'lutff_1/cout')

wire n151;
// (1, 5, 'lutff_3/cout')

wire n152;
// (6, 3, 'lutff_4/cout')

wire n153;
// (1, 4, 'lutff_1/cout')

wire n154;
// (1, 3, 'lutff_5/cout')

wire n155;
// (6, 4, 'lutff_2/cout')

wire n156;
// (1, 1, 'lutff_5/cout')

wire n157;
// (5, 3, 'lutff_1/cout')

wire n158;
// (7, 3, 'lutff_3/cout')

wire n159;
// (1, 5, 'lutff_5/cout')

wire n160;
// (6, 3, 'lutff_6/cout')

wire n161;
// (5, 3, 'lutff_3/lout')

wire n162;
// (5, 4, 'lutff_2/out')

wire n163;
// (5, 4, 'lutff_2/lout')

wire n164;
// (7, 3, 'lutff_5/out')

wire n165;
// (7, 3, 'lutff_5/lout')

wire n166;
// (1, 5, 'lutff_7/lout')

wire n167;
// (1, 3, 'lutff_0/out')

wire n168;
// (1, 3, 'lutff_0/lout')

wire n169;
// (1, 3, 'carry_in_mux')

// Carry-In for (1 3)
assign n169 = 1;

wire n170;
// (5, 5, 'lutff_3/lout')

wire n171;
// (2, 4, 'lutff_5/lout')

wire n172;
// (1, 1, 'lutff_0/out')

wire n173;
// (1, 1, 'lutff_0/lout')

wire n174;
// (1, 1, 'carry_in_mux')

// Carry-In for (1 1)
assign n174 = 1;

wire n175;
// (5, 3, 'lutff_5/out')

wire n176;
// (5, 3, 'lutff_5/lout')

wire n177;
// (5, 4, 'lutff_4/lout')

wire n178;
// (1, 5, 'lutff_0/out')

wire n179;
// (1, 5, 'lutff_0/lout')

wire n180;
// (1, 5, 'carry_in_mux')

// Carry-In for (1 5)
assign n180 = 1;

wire n181;
// (7, 3, 'lutff_7/out')

wire n182;
// (7, 3, 'lutff_7/lout')

wire n183;
// (4, 4, 'lutff_3/lout')

wire n184;
// (1, 3, 'lutff_2/lout')

wire n185;
// (4, 3, 'lutff_1/out')

wire n186;
// (4, 3, 'lutff_1/lout')

wire n187;
// (2, 4, 'lutff_7/lout')

wire n188;
// (1, 1, 'lutff_2/out')

wire n189;
// (1, 1, 'lutff_2/lout')

wire n190;
// (7, 3, 'lutff_0/out')

wire n191;
// (7, 3, 'lutff_0/lout')

wire n192;
// (7, 3, 'carry_in_mux')

// Carry-In for (7 3)
assign n192 = 1;

wire n193;
// (5, 3, 'lutff_7/out')

wire n194;
// (5, 3, 'lutff_7/lout')

wire n195;
// (5, 4, 'lutff_6/lout')

wire n196;
// (1, 5, 'lutff_2/out')

wire n197;
// (1, 5, 'lutff_2/lout')

wire n198;
// (4, 4, 'lutff_5/lout')

wire n199;
// (1, 3, 'lutff_4/lout')

wire n200;
// (5, 5, 'lutff_7/lout')

wire n201;
// (1, 4, 'lutff_3/lout')

wire n202;
// (2, 4, 'lutff_0/lout')

wire n203;
// (1, 1, 'lutff_4/out')

wire n204;
// (1, 1, 'lutff_4/lout')

wire n205;
// (5, 3, 'lutff_0/out')

wire n206;
// (5, 3, 'lutff_0/lout')

wire n207;
// (5, 3, 'carry_in_mux')

// Carry-In for (5 3)
assign n207 = 1;

wire n208;
// (7, 3, 'lutff_2/out')

wire n209;
// (7, 3, 'lutff_2/lout')

wire n210;
// (7, 4, 'lutff_1/lout')

wire n211;
// (1, 5, 'lutff_4/lout')

wire n212;
// (4, 4, 'lutff_7/lout')

wire n213;
// (1, 3, 'lutff_6/lout')

wire n214;
// (1, 4, 'lutff_5/lout')

wire n215;
// (2, 4, 'lutff_2/lout')

wire n216;
// (2, 3, 'lutff_6/lout')

wire n217;
// (5, 3, 'lutff_2/lout')

wire n218;
// (5, 4, 'lutff_1/out')

wire n219;
// (5, 4, 'lutff_1/lout')

wire n220;
// (7, 3, 'lutff_4/out')

wire n221;
// (7, 3, 'lutff_4/lout')

wire n222;
// (1, 5, 'lutff_6/out')

wire n223;
// (1, 5, 'lutff_6/lout')

wire n224;
// (6, 3, 'lutff_1/out')

wire n225;
// (6, 3, 'lutff_1/lout')

wire n226;
// (4, 4, 'lutff_0/lout')

wire n227;
// (1, 2, 'lutff_1/out')

wire n228;
// (1, 2, 'lutff_1/lout')

wire n229;
// (1, 4, 'lutff_7/lout')

wire n230;
// (4, 3, 'lutff_6/lout')

wire n231;
// (5, 4, 'lutff_3/out')

wire n232;
// (5, 4, 'lutff_3/lout')

wire n233;
// (6, 3, 'lutff_3/out')

wire n234;
// (6, 3, 'lutff_3/lout')

wire n235;
// (4, 4, 'lutff_2/lout')

wire n236;
// (1, 3, 'lutff_1/lout')

wire n237;
// (1, 2, 'lutff_3/out')

wire n238;
// (1, 2, 'lutff_3/lout')

wire n239;
// (1, 4, 'lutff_0/lout')

wire n240;
// (2, 3, 'lutff_1/out')

wire n241;
// (2, 3, 'lutff_1/lout')

wire n242;
// (4, 3, 'lutff_3/lout')

wire n243;
// (6, 4, 'lutff_1/lout')

wire n244;
// (5, 4, 'lutff_5/lout')

wire n245;
// (1, 5, 'lutff_1/out')

wire n246;
// (1, 5, 'lutff_1/lout')

wire n247;
// (6, 3, 'lutff_5/out')

wire n248;
// (6, 3, 'lutff_5/lout')

wire n249;
// (1, 3, 'lutff_3/lout')

wire n250;
// (1, 4, 'lutff_2/lout')

wire n251;
// (2, 3, 'lutff_3/lout')

wire n252;
// (4, 3, 'lutff_5/lout')

wire n253;
// (6, 4, 'lutff_3/out')

wire n254;
// (6, 4, 'lutff_3/lout')

wire n255;
// (7, 4, 'lutff_0/lout')

wire n256;
// (1, 1, 'lutff_6/out')

wire n257;
// (1, 1, 'lutff_6/lout')

wire n258;
// (6, 3, 'lutff_7/lout')

wire n259;
// (4, 4, 'lutff_6/lout')

wire n260;
// (4, 5, 'lutff_5/lout')

wire n261;
// (1, 4, 'lutff_4/lout')

wire n262;
// (2, 3, 'lutff_5/lout')

wire n263;
// (2, 4, 'lutff_4/lout')

wire n264;
// (4, 3, 'lutff_7/lout')

wire n265;
// (6, 4, 'lutff_5/lout')

wire n266;
// (5, 4, 'lutff_0/out')

wire n267;
// (5, 4, 'lutff_0/lout')

wire n268;
// (7, 4, 'lutff_2/lout')

wire n269;
// (5, 3, 'lutff_4/out')

wire n270;
// (5, 3, 'lutff_4/lout')

wire n271;
// (7, 3, 'lutff_6/out')

wire n272;
// (7, 3, 'lutff_6/lout')

wire n273;
// (6, 3, 'lutff_0/out')

wire n274;
// (6, 3, 'lutff_0/lout')

wire n275;
// (6, 3, 'carry_in_mux')

// Carry-In for (6 3)
assign n275 = 1;

wire n276;
// (2, 5, 'lutff_5/lout')

wire n277;
// (1, 2, 'lutff_0/out')

wire n278;
// (1, 2, 'lutff_0/lout')

wire n279;
// (1, 4, 'lutff_6/lout')

wire n280;
// (5, 5, 'lutff_4/lout')

wire n281;
// (4, 3, 'lutff_0/out')

wire n282;
// (4, 3, 'lutff_0/lout')

wire n283;
// (4, 3, 'carry_in_mux')

// Carry-In for (4 3)
assign n283 = 1;

wire n284;
// (2, 3, 'lutff_7/lout')

wire n285;
// (2, 4, 'lutff_6/lout')

wire n286;
// (6, 4, 'lutff_7/lout')

wire n287;
// (1, 1, 'lutff_1/out')

wire n288;
// (1, 1, 'lutff_1/lout')

wire n289;
// (5, 3, 'lutff_6/out')

wire n290;
// (5, 3, 'lutff_6/lout')

wire n291;
// (6, 3, 'lutff_2/out')

wire n292;
// (6, 3, 'lutff_2/lout')

wire n293;
// (4, 4, 'lutff_1/lout')

wire n294;
// (2, 5, 'lutff_7/lout')

wire n295;
// (1, 2, 'lutff_2/out')

wire n296;
// (1, 2, 'lutff_2/lout')

wire n297;
// (2, 3, 'lutff_0/out')

wire n298;
// (2, 3, 'lutff_0/lout')

wire n299;
// (2, 3, 'carry_in_mux')

// Carry-In for (2 3)
assign n299 = 1;

wire n300;
// (6, 4, 'lutff_0/lout')

wire n301;
// (4, 3, 'lutff_2/lout')

wire n302;
// (1, 1, 'lutff_3/out')

wire n303;
// (1, 1, 'lutff_3/lout')

wire n304;
// (7, 3, 'lutff_1/out')

wire n305;
// (7, 3, 'lutff_1/lout')

wire n306;
// (5, 4, 'lutff_7/lout')

wire n307;
// (1, 5, 'lutff_3/out')

wire n308;
// (1, 5, 'lutff_3/lout')

wire n309;
// (2, 5, 'lutff_0/lout')

wire n310;
// (6, 3, 'lutff_4/lout')

wire n311;
// (1, 2, 'lutff_4/lout')

wire n312;
// (1, 4, 'lutff_1/lout')

wire n313;
// (1, 3, 'lutff_5/lout')

wire n314;
// (2, 3, 'lutff_2/lout')

wire n315;
// (2, 4, 'lutff_1/lout')

wire n316;
// (4, 3, 'lutff_4/lout')

wire n317;
// (6, 4, 'lutff_2/out')

wire n318;
// (6, 4, 'lutff_2/lout')

wire n319;
// (1, 1, 'lutff_5/out')

wire n320;
// (1, 1, 'lutff_5/lout')

wire n321;
// (5, 3, 'lutff_1/lout')

wire n322;
// (7, 3, 'lutff_3/lout')

wire n323;
// (1, 5, 'lutff_5/out')

wire n324;
// (1, 5, 'lutff_5/lout')

wire n325;
// (6, 3, 'lutff_6/lout')

wire n326;
// (1, 3, 'lutff_7/lout')

wire n327;
// (2, 3, 'lutff_4/lout')

wire n328;
// (2, 4, 'lutff_3/lout')

wire n329;
// (6, 4, 'lutff_4/lout')

wire n330;
// (1, 1, 'lutff_7/out')

wire n331;
// (1, 1, 'lutff_7/lout')

assign n163 = /* LUT    5  4  2 */ 1'b0;
assign n165 = /* LUT    7  3  5 */ 1'b0;
assign n168 = /* LUT    1  3  0 */ 1'b0;
assign n173 = /* LUT    1  1  0 */ 1'b0;
assign n176 = /* LUT    5  3  5 */ 1'b0;
assign n179 = /* LUT    1  5  0 */ 1'b0;
assign n182 = /* LUT    7  3  7 */ 1'b0;
assign n186 = /* LUT    4  3  1 */ 1'b0;
assign n189 = /* LUT    1  1  2 */ 1'b0;
assign n191 = /* LUT    7  3  0 */ 1'b0;
assign n194 = /* LUT    5  3  7 */ 1'b0;
assign n197 = /* LUT    1  5  2 */ 1'b0;
assign n204 = /* LUT    1  1  4 */ 1'b0;
assign n206 = /* LUT    5  3  0 */ 1'b0;
assign n209 = /* LUT    7  3  2 */ 1'b0;
assign n219 = /* LUT    5  4  1 */ 1'b0;
assign n221 = /* LUT    7  3  4 */ 1'b0;
assign n223 = /* LUT    1  5  6 */ 1'b0;
assign n225 = /* LUT    6  3  1 */ 1'b0;
assign n228 = /* LUT    1  2  1 */ 1'b0;
assign n232 = /* LUT    5  4  3 */ 1'b0;
assign n234 = /* LUT    6  3  3 */ 1'b0;
assign n238 = /* LUT    1  2  3 */ 1'b0;
assign n241 = /* LUT    2  3  1 */ 1'b0;
assign n246 = /* LUT    1  5  1 */ 1'b0;
assign n248 = /* LUT    6  3  5 */ 1'b0;
assign n254 = /* LUT    6  4  3 */ 1'b0;
assign n257 = /* LUT    1  1  6 */ 1'b0;
assign n267 = /* LUT    5  4  0 */ 1'b0;
assign n270 = /* LUT    5  3  4 */ 1'b0;
assign n272 = /* LUT    7  3  6 */ 1'b0;
assign n274 = /* LUT    6  3  0 */ 1'b0;
assign n278 = /* LUT    1  2  0 */ 1'b0;
assign n282 = /* LUT    4  3  0 */ 1'b0;
assign n288 = /* LUT    1  1  1 */ 1'b0;
assign n290 = /* LUT    5  3  6 */ 1'b0;
assign n292 = /* LUT    6  3  2 */ 1'b0;
assign n296 = /* LUT    1  2  2 */ 1'b0;
assign n298 = /* LUT    2  3  0 */ 1'b0;
assign n303 = /* LUT    1  1  3 */ 1'b0;
assign n305 = /* LUT    7  3  1 */ 1'b0;
assign n308 = /* LUT    1  5  3 */ 1'b0;
assign n318 = /* LUT    6  4  2 */ 1'b0;
assign n320 = /* LUT    1  1  5 */ 1'b0;
assign n324 = /* LUT    1  5  5 */ 1'b0;
assign n331 = /* LUT    1  1  7 */ 1'b0;
assign n161 = /* LUT    5  3  3 */ !n57;
assign n166 = /* LUT    1  5  7 */ (n43 ? (n42 ? (n17 ? n38 : 1'b0) : 1'b0) : 1'b1);
assign n170 = /* LUT    5  5  3 */ (n80 ? (n81 ? (n87 ? 1'b0 : n95) : n95) : n95);
assign n171 = /* LUT    2  4  5 */ (n30 ? 1'b0 : (n32 ? 1'b0 : (n29 ? 1'b0 : !n28)));
assign n177 = /* LUT    5  4  4 */ (n99 ? (n96 ? (n66 ? n64 : 1'b0) : 1'b0) : 1'b1);
assign n183 = /* LUT    4  4  3 */ (n85 ? !n63 : n63);
assign n184 = /* LUT    1  3  2 */ !n28;
assign n187 = /* LUT    2  4  7 */ (n16 ? 1'b0 : (n31 ? 1'b0 : (n36 ? 1'b0 : !n34)));
assign n195 = /* LUT    5  4  6 */ (n59 ? (n51 ? 1'b0 : (n60 ? n58 : 1'b0)) : 1'b0);
assign n198 = /* LUT    4  4  5 */ (n65 ? 1'b0 : (n71 ? 1'b0 : (n57 ? n56 : 1'b0)));
assign n199 = /* LUT    1  3  4 */ !n30;
assign n200 = /* LUT    5  5  7 */ (n63 ? 1'b0 : (n71 ? 1'b0 : (n62 ? 1'b0 : !n65)));
assign n201 = /* LUT    1  4  3 */ !n36;
assign n202 = /* LUT    2  4  0 */ (n50 ? !n34 : n34);
assign n210 = /* LUT    7  4  1 */ !n63;
assign n211 = /* LUT    1  5  4 */ !n21;
assign n212 = /* LUT    4  4  7 */ (n60 ? 1'b0 : (n61 ? (n62 ? 1'b0 : !n63) : 1'b0));
assign n213 = /* LUT    1  3  6 */ !n25;
assign n214 = /* LUT    1  4  5 */ !n16;
assign n215 = /* LUT    2  4  2 */ (n54 ? !n35 : n35);
assign n216 = /* LUT    2  3  6 */ (n48 ? !n25 : n25);
assign n217 = /* LUT    5  3  2 */ !n56;
assign n226 = /* LUT    4  4  0 */ (n79 ? !n60 : n60);
assign n229 = /* LUT    1  4  7 */ (n16 ? (n34 ? (n32 ? n28 : 1'b0) : 1'b0) : 1'b0);
assign n230 = /* LUT    4  3  6 */ (n77 ? !n58 : n58);
assign n235 = /* LUT    4  4  2 */ (n84 ? !n62 : n62);
assign n236 = /* LUT    1  3  1 */ !n32;
assign n239 = /* LUT    1  4  0 */ !n34;
assign n242 = /* LUT    4  3  3 */ (n74 ? !n57 : n57);
assign n243 = /* LUT    6  4  1 */ !n61;
assign n244 = /* LUT    5  4  5 */ (n71 ? (n56 ? 1'b0 : (n57 ? n65 : 1'b0)) : 1'b0);
assign n249 = /* LUT    1  3  3 */ !n29;
assign n250 = /* LUT    1  4  2 */ !n35;
assign n251 = /* LUT    2  3  3 */ (n45 ? !n29 : n29);
assign n252 = /* LUT    4  3  5 */ (n76 ? !n52 : n52);
assign n255 = /* LUT    7  4  0 */ !n62;
assign n258 = /* LUT    6  3  7 */ !n59;
assign n259 = /* LUT    4  4  6 */ (n71 ? !n65 : n65);
assign n260 = /* LUT    4  5  5 */ (n25 ? n86 : (n86 ? (n26 ? !n24 : 1'b1) : 1'b0));
assign n261 = /* LUT    1  4  4 */ n40;
assign n262 = /* LUT    2  3  5 */ (n47 ? !n31 : n31);
assign n263 = /* LUT    2  4  4 */ (n32 ? !n16 : n16);
assign n264 = /* LUT    4  3  7 */ (n78 ? !n59 : n59);
assign n265 = /* LUT    6  4  5 */ !n71;
assign n268 = /* LUT    7  4  2 */ (n103 ? (n66 ? (n96 ? !n67 : 1'b1) : 1'b1) : 1'b0);
assign n276 = /* LUT    2  5  5 */ n19;
assign n279 = /* LUT    1  4  6 */ n15;
assign n280 = /* LUT    5  5  4 */ n91;
assign n284 = /* LUT    2  3  7 */ (n49 ? !n26 : n26);
assign n285 = /* LUT    2  4  6 */ (n30 ? (n36 ? 1'b0 : (n31 ? 1'b0 : n29)) : 1'b0);
assign n286 = /* LUT    6  4  7 */ (n59 ? 1'b0 : (n52 ? 1'b0 : (n58 ? 1'b0 : !n51)));
assign n293 = /* LUT    4  4  1 */ (n83 ? !n61 : n61);
assign n294 = /* LUT    2  5  7 */ (n25 ? 1'b0 : (n35 ? 1'b0 : (n21 ? !n26 : 1'b0)));
assign n300 = /* LUT    6  4  0 */ !n60;
assign n301 = /* LUT    4  3  2 */ (n73 ? !n56 : n56);
assign n306 = /* LUT    5  4  7 */ (n61 ? 1'b0 : (n57 ? 1'b0 : (n52 ? !n56 : 1'b0)));
assign n309 = /* LUT    2  5  0 */ (n35 ? 1'b0 : (n37 ? (n39 ? n21 : 1'b0) : 1'b0));
assign n310 = /* LUT    6  3  4 */ !n51;
assign n311 = /* LUT    1  2  4 */ (n27 ? (n25 ? (n24 ? !n26 : 1'b1) : 1'b1) : 1'b0);
assign n312 = /* LUT    1  4  1 */ 1'b1;
assign n313 = /* LUT    1  3  5 */ !n31;
assign n314 = /* LUT    2  3  2 */ (n44 ? !n28 : n28);
assign n315 = /* LUT    2  4  1 */ (n53 ? !n21 : n21);
assign n316 = /* LUT    4  3  4 */ (n75 ? !n51 : n51);
assign n321 = /* LUT    5  3  1 */ !n65;
assign n322 = /* LUT    7  3  3 */ !n52;
assign n325 = /* LUT    6  3  6 */ !n58;
assign n326 = /* LUT    1  3  7 */ !n26;
assign n327 = /* LUT    2  3  4 */ (n46 ? !n30 : n30);
assign n328 = /* LUT    2  4  3 */ (n55 ? !n36 : n36);
assign n329 = /* LUT    6  4  4 */ (n101 ? n14 : 1'b0);
assign n104 = /* CARRY  5  3  3 */ (n11 & n70) | ((n11 | n70) & n121);
assign n105 = /* CARRY  5  4  2 */ (1'b0 & n97) | ((1'b0 | n97) & n122);
assign n106 = /* CARRY  7  3  5 */ (n90 & 1'b0) | ((n90 | 1'b0) & n123);
assign n107 = /* CARRY  1  3  0 */ (1'b0 & n15) | ((1'b0 | n15) & n169);
assign n108 = /* CARRY  1  1  0 */ (1'b0 & n15) | ((1'b0 | n15) & n174);
assign n109 = /* CARRY  5  3  5 */ (1'b0 & n82) | ((1'b0 | n82) & n138);
assign n110 = /* CARRY  1  5  0 */ (n7 & 1'b0) | ((n7 | 1'b0) & n180);
assign n102 = /* CARRY  7  3  7 */ (n94 & n11) | ((n94 | n11) & n139);
assign n111 = /* CARRY  1  3  2 */ (1'b0 & n4) | ((1'b0 | n4) & n127);
assign n73  = /* CARRY  4  3  1 */ (n65 & 1'b0) | ((n65 | 1'b0) & n142);
assign n112 = /* CARRY  1  1  2 */ (1'b0 & n4) | ((1'b0 | n4) & n143);
assign n113 = /* CARRY  7  3  0 */ (n69 & 1'b0) | ((n69 | 1'b0) & n192);
assign n92  = /* CARRY  5  3  7 */ (n90 & 1'b0) | ((n90 | 1'b0) & n144);
assign n114 = /* CARRY  1  5  2 */ (1'b0 & n9) | ((1'b0 | n9) & n130);
assign n115 = /* CARRY  1  3  4 */ (n6 & 1'b0) | ((n6 | 1'b0) & n132);
assign n40  = /* CARRY  1  4  3 */ (1'b0 & n13) | ((1'b0 | n13) & n133);
assign n53  = /* CARRY  2  4  0 */ (n34 & 1'b0) | ((n34 | 1'b0) & n50);
assign n116 = /* CARRY  1  1  4 */ (n6 & 1'b0) | ((n6 | 1'b0) & n149);
assign n117 = /* CARRY  5  3  0 */ (n91 & 1'b0) | ((n91 | 1'b0) & n207);
assign n118 = /* CARRY  7  3  2 */ (1'b0 & n88) | ((1'b0 | n88) & n150);
assign n103 = /* CARRY  7  4  1 */ (1'b0 & n98) | ((1'b0 | n98) & n134);
assign n119 = /* CARRY  1  5  4 */ (n11 & n18) | ((n11 | n18) & n151);
assign n120 = /* CARRY  1  3  6 */ (1'b0 & n8) | ((1'b0 | n8) & n154);
assign n55  = /* CARRY  2  4  2 */ (1'b0 & n35) | ((1'b0 | n35) & n54);
assign n49  = /* CARRY  2  3  6 */ (n25 & 1'b0) | ((n25 | 1'b0) & n48);
assign n121 = /* CARRY  5  3  2 */ (n11 & n69) | ((n11 | n69) & n157);
assign n122 = /* CARRY  5  4  1 */ (n11 & n94) | ((n11 | n94) & n137);
assign n123 = /* CARRY  7  3  4 */ (n89 & 1'b0) | ((n89 | 1'b0) & n158);
assign n43  = /* CARRY  1  5  6 */ (1'b0 & n13) | ((1'b0 | n13) & n159);
assign n124 = /* CARRY  6  3  1 */ (n68 & 1'b0) | ((n68 | 1'b0) & n140);
assign n83  = /* CARRY  4  4  0 */ (1'b0 & n60) | ((1'b0 | n60) & n79);
assign n125 = /* CARRY  1  2  1 */ (n18 & n11) | ((n18 | n11) & n141);
assign n78  = /* CARRY  4  3  6 */ (n58 & 1'b0) | ((n58 | 1'b0) & n77);
assign n99  = /* CARRY  5  4  3 */ (1'b0 & n98) | ((1'b0 | n98) & n105);
assign n126 = /* CARRY  6  3  3 */ (n70 & 1'b0) | ((n70 | 1'b0) & n145);
assign n85  = /* CARRY  4  4  2 */ (1'b0 & n62) | ((1'b0 | n62) & n84);
assign n127 = /* CARRY  1  3  1 */ (n3 & 1'b0) | ((n3 | 1'b0) & n107);
assign n27  = /* CARRY  1  2  3 */ (1'b0 & n13) | ((1'b0 | n13) & n146);
assign n128 = /* CARRY  1  4  0 */ (1'b0 & n10) | ((1'b0 | n10) & n33);
assign n44  = /* CARRY  2  3  1 */ (n32 & 1'b0) | ((n32 | 1'b0) & n147);
assign n75  = /* CARRY  4  3  3 */ (n57 & 1'b0) | ((n57 | 1'b0) & n74);
assign n129 = /* CARRY  6  4  1 */ (1'b0 & n94) | ((1'b0 | n94) & n148);
assign n130 = /* CARRY  1  5  1 */ (n8 & 1'b0) | ((n8 | 1'b0) & n110);
assign n131 = /* CARRY  6  3  5 */ (n11 & n82) | ((n11 | n82) & n152);
assign n132 = /* CARRY  1  3  3 */ (n5 & 1'b0) | ((n5 | 1'b0) & n111);
assign n133 = /* CARRY  1  4  2 */ (1'b0 & n12) | ((1'b0 | n12) & n153);
assign n46  = /* CARRY  2  3  3 */ (1'b0 & n29) | ((1'b0 | n29) & n45);
assign n77  = /* CARRY  4  3  5 */ (n52 & 1'b0) | ((n52 | 1'b0) & n76);
assign n101 = /* CARRY  6  4  3 */ (1'b0 & n98) | ((1'b0 | n98) & n155);
assign n134 = /* CARRY  7  4  0 */ (n97 & 1'b0) | ((n97 | 1'b0) & n102);
assign n135 = /* CARRY  1  1  6 */ (n8 & n11) | ((n8 | n11) & n156);
assign n100 = /* CARRY  6  3  7 */ (n11 & n90) | ((n11 | n90) & n160);
assign n136 = /* CARRY  1  4  4 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n40);
assign n48  = /* CARRY  2  3  5 */ (n31 & 1'b0) | ((n31 | 1'b0) & n47);
assign n79  = /* CARRY  4  3  7 */ (n59 & 1'b0) | ((n59 | 1'b0) & n78);
assign n137 = /* CARRY  5  4  0 */ (n93 & 1'b0) | ((n93 | 1'b0) & n92);
assign n138 = /* CARRY  5  3  4 */ (1'b0 & n88) | ((1'b0 | n88) & n104);
assign n139 = /* CARRY  7  3  6 */ (1'b0 & n93) | ((1'b0 | n93) & n106);
assign n140 = /* CARRY  6  3  0 */ (n91 & 1'b0) | ((n91 | 1'b0) & n275);
assign n141 = /* CARRY  1  2  0 */ (1'b0 & n10) | ((1'b0 | n10) & n22);
assign n142 = /* CARRY  4  3  0 */ (1'b0 & n71) | ((1'b0 | n71) & n283);
assign n50  = /* CARRY  2  3  7 */ (1'b0 & n26) | ((1'b0 | n26) & n49);
assign n143 = /* CARRY  1  1  1 */ (1'b0 & n3) | ((1'b0 | n3) & n108);
assign n144 = /* CARRY  5  3  6 */ (n89 & 1'b0) | ((n89 | 1'b0) & n109);
assign n145 = /* CARRY  6  3  2 */ (n69 & 1'b0) | ((n69 | 1'b0) & n124);
assign n84  = /* CARRY  4  4  1 */ (1'b0 & n61) | ((1'b0 | n61) & n83);
assign n146 = /* CARRY  1  2  2 */ (n12 & 1'b0) | ((n12 | 1'b0) & n125);
assign n147 = /* CARRY  2  3  0 */ (1'b0 & n16) | ((1'b0 | n16) & n299);
assign n148 = /* CARRY  6  4  0 */ (n11 & n93) | ((n11 | n93) & n100);
assign n74  = /* CARRY  4  3  2 */ (1'b0 & n56) | ((1'b0 | n56) & n73);
assign n149 = /* CARRY  1  1  3 */ (n5 & 1'b0) | ((n5 | 1'b0) & n112);
assign n150 = /* CARRY  7  3  1 */ (n70 & n11) | ((n70 | n11) & n113);
assign n151 = /* CARRY  1  5  3 */ (n11 & n10) | ((n11 | n10) & n114);
assign n152 = /* CARRY  6  3  4 */ (n88 & 1'b0) | ((n88 | 1'b0) & n126);
assign n153 = /* CARRY  1  4  1 */ (n11 & n18) | ((n11 | n18) & n128);
assign n154 = /* CARRY  1  3  5 */ (1'b0 & n7) | ((1'b0 | n7) & n115);
assign n45  = /* CARRY  2  3  2 */ (1'b0 & n28) | ((1'b0 | n28) & n44);
assign n54  = /* CARRY  2  4  1 */ (1'b0 & n21) | ((1'b0 | n21) & n53);
assign n76  = /* CARRY  4  3  4 */ (n51 & 1'b0) | ((n51 | 1'b0) & n75);
assign n155 = /* CARRY  6  4  2 */ (1'b0 & n97) | ((1'b0 | n97) & n129);
assign n156 = /* CARRY  1  1  5 */ (n7 & 1'b0) | ((n7 | 1'b0) & n116);
assign n157 = /* CARRY  5  3  1 */ (1'b0 & n68) | ((1'b0 | n68) & n117);
assign n158 = /* CARRY  7  3  3 */ (1'b0 & n82) | ((1'b0 | n82) & n118);
assign n159 = /* CARRY  1  5  5 */ (n12 & 1'b0) | ((n12 | 1'b0) & n119);
assign n160 = /* CARRY  6  3  6 */ (n89 & n11) | ((n89 | n11) & n131);
assign n33  = /* CARRY  1  3  7 */ (n9 & n11) | ((n9 | n11) & n120);
assign n47  = /* CARRY  2  3  4 */ (1'b0 & n30) | ((1'b0 | n30) & n46);
assign n22  = /* CARRY  1  1  7 */ (n11 & n9) | ((n11 | n9) & n135);
/* FF  5  3  3 */ assign n70 = n161;
/* FF  5  4  2 */ assign n162 = n163;
/* FF  7  3  5 */ assign n164 = n165;
/* FF  1  5  7 */ assign n19 = n166;
/* FF  1  3  0 */ assign n167 = n168;
/* FF  5  5  3 */ assign n86 = n170;
/* FF  2  4  5 */ assign n37 = n171;
/* FF  1  1  0 */ assign n172 = n173;
/* FF  5  3  5 */ assign n175 = n176;
/* FF  5  4  4 */ assign n72 = n177;
/* FF  1  5  0 */ assign n178 = n179;
/* FF  7  3  7 */ assign n181 = n182;
/* FF  4  4  3 */ always @(posedge io_0_8_1) if (n19) n63 <= n72 ? 1'b0 : n183;
/* FF  1  3  2 */ assign n4 = n184;
/* FF  4  3  1 */ assign n185 = n186;
/* FF  2  4  7 */ assign n39 = n187;
/* FF  1  1  2 */ assign n188 = n189;
/* FF  7  3  0 */ assign n190 = n191;
/* FF  5  3  7 */ assign n193 = n194;
/* FF  5  4  6 */ assign n80 = n195;
/* FF  1  5  2 */ assign n196 = n197;
/* FF  4  4  5 */ assign n64 = n198;
/* FF  1  3  4 */ assign n6 = n199;
/* FF  5  5  7 */ assign n87 = n200;
/* FF  1  4  3 */ assign n13 = n201;
/* FF  2  4  0 */ always @(posedge io_0_8_1) if (1'b1) n34 <= n41 ? 1'b0 : n202;
/* FF  1  1  4 */ assign n203 = n204;
/* FF  5  3  0 */ assign n205 = n206;
/* FF  7  3  2 */ assign n208 = n209;
/* FF  7  4  1 */ assign n98 = n210;
/* FF  1  5  4 */ assign n18 = n211;
/* FF  4  4  7 */ assign n66 = n212;
/* FF  1  3  6 */ assign n8 = n213;
/* FF  1  4  5 */ assign n15 = n214;
/* FF  2  4  2 */ always @(posedge io_0_8_1) if (1'b1) n35 <= n41 ? 1'b0 : n215;
/* FF  2  3  6 */ always @(posedge io_0_8_1) if (1'b1) n25 <= n19 ? 1'b0 : n216;
/* FF  5  3  2 */ assign n69 = n217;
/* FF  5  4  1 */ assign n218 = n219;
/* FF  7  3  4 */ assign n220 = n221;
/* FF  1  5  6 */ assign n222 = n223;
/* FF  6  3  1 */ assign n224 = n225;
/* FF  4  4  0 */ always @(posedge io_0_8_1) if (n19) n60 <= n72 ? 1'b0 : n226;
/* FF  1  2  1 */ assign n227 = n228;
/* FF  1  4  7 */ assign n17 = n229;
/* FF  4  3  6 */ always @(posedge io_0_8_1) if (n19) n58 <= n72 ? 1'b0 : n230;
/* FF  5  4  3 */ assign n231 = n232;
/* FF  6  3  3 */ assign n233 = n234;
/* FF  4  4  2 */ always @(posedge io_0_8_1) if (n19) n62 <= n72 ? 1'b0 : n235;
/* FF  1  3  1 */ assign n3 = n236;
/* FF  1  2  3 */ assign n237 = n238;
/* FF  1  4  0 */ assign n10 = n239;
/* FF  2  3  1 */ assign n240 = n241;
/* FF  4  3  3 */ always @(posedge io_0_8_1) if (n19) n57 <= n72 ? 1'b0 : n242;
/* FF  6  4  1 */ assign n94 = n243;
/* FF  5  4  5 */ assign n67 = n244;
/* FF  1  5  1 */ assign n245 = n246;
/* FF  6  3  5 */ assign n247 = n248;
/* FF  1  3  3 */ assign n5 = n249;
/* FF  1  4  2 */ assign n12 = n250;
/* FF  2  3  3 */ always @(posedge io_0_8_1) if (1'b1) n29 <= n19 ? 1'b0 : n251;
/* FF  4  3  5 */ always @(posedge io_0_8_1) if (n19) n52 <= n72 ? 1'b0 : n252;
/* FF  6  4  3 */ assign n253 = n254;
/* FF  7  4  0 */ assign n97 = n255;
/* FF  1  1  6 */ assign n256 = n257;
/* FF  6  3  7 */ assign n90 = n258;
/* FF  4  4  6 */ always @(posedge io_0_8_1) if (n19) n65 <= n72 ? 1'b0 : n259;
/* FF  4  5  5 */ always @(posedge io_0_8_1) if (1'b1) io_3_0_0 <= 1'b0 ? 1'b0 : n260;
/* FF  1  4  4 */ assign n14 = n261;
/* FF  2  3  5 */ always @(posedge io_0_8_1) if (1'b1) n31 <= n19 ? 1'b0 : n262;
/* FF  2  4  4 */ always @(posedge io_0_8_1) if (1'b1) n32 <= n41 ? 1'b0 : n263;
/* FF  4  3  7 */ always @(posedge io_0_8_1) if (n19) n59 <= n72 ? 1'b0 : n264;
/* FF  6  4  5 */ assign n91 = n265;
/* FF  5  4  0 */ assign n266 = n267;
/* FF  7  4  2 */ always @(posedge io_0_8_1) if (1'b1) io_2_0_1 <= 1'b0 ? 1'b0 : n268;
/* FF  5  3  4 */ assign n269 = n270;
/* FF  7  3  6 */ assign n271 = n272;
/* FF  6  3  0 */ assign n273 = n274;
/* FF  2  5  5 */ assign n41 = n276;
/* FF  1  2  0 */ assign n277 = n278;
/* FF  1  4  6 */ always @(posedge io_0_8_1) if (1'b1) n16 <= n19 ? 1'b0 : n279;
/* FF  5  5  4 */ always @(posedge io_0_8_1) if (n19) n71 <= n72 ? 1'b0 : n280;
/* FF  4  3  0 */ assign n281 = n282;
/* FF  2  3  7 */ always @(posedge io_0_8_1) if (1'b1) n26 <= n19 ? 1'b0 : n284;
/* FF  2  4  6 */ assign n38 = n285;
/* FF  6  4  7 */ assign n96 = n286;
/* FF  1  1  1 */ assign n287 = n288;
/* FF  5  3  6 */ assign n289 = n290;
/* FF  6  3  2 */ assign n291 = n292;
/* FF  4  4  1 */ always @(posedge io_0_8_1) if (n19) n61 <= n72 ? 1'b0 : n293;
/* FF  2  5  7 */ assign n42 = n294;
/* FF  1  2  2 */ assign n295 = n296;
/* FF  2  3  0 */ assign n297 = n298;
/* FF  6  4  0 */ assign n93 = n300;
/* FF  4  3  2 */ always @(posedge io_0_8_1) if (n19) n56 <= n72 ? 1'b0 : n301;
/* FF  1  1  3 */ assign n302 = n303;
/* FF  7  3  1 */ assign n304 = n305;
/* FF  5  4  7 */ assign n81 = n306;
/* FF  1  5  3 */ assign n307 = n308;
/* FF  2  5  0 */ assign n24 = n309;
/* FF  6  3  4 */ assign n88 = n310;
/* FF  1  2  4 */ always @(posedge io_0_8_1) if (1'b1) io_2_0_0 <= 1'b0 ? 1'b0 : n311;
/* FF  1  4  1 */ assign n11 = n312;
/* FF  1  3  5 */ assign n7 = n313;
/* FF  2  3  2 */ always @(posedge io_0_8_1) if (1'b1) n28 <= n19 ? 1'b0 : n314;
/* FF  2  4  1 */ always @(posedge io_0_8_1) if (1'b1) n21 <= n41 ? 1'b0 : n315;
/* FF  4  3  4 */ always @(posedge io_0_8_1) if (n19) n51 <= n72 ? 1'b0 : n316;
/* FF  6  4  2 */ assign n317 = n318;
/* FF  1  1  5 */ assign n319 = n320;
/* FF  5  3  1 */ assign n68 = n321;
/* FF  7  3  3 */ assign n82 = n322;
/* FF  1  5  5 */ assign n323 = n324;
/* FF  6  3  6 */ assign n89 = n325;
/* FF  1  3  7 */ assign n9 = n326;
/* FF  2  3  4 */ always @(posedge io_0_8_1) if (1'b1) n30 <= n19 ? 1'b0 : n327;
/* FF  2  4  3 */ always @(posedge io_0_8_1) if (1'b1) n36 <= n41 ? 1'b0 : n328;
/* FF  6  4  4 */ assign n95 = n329;
/* FF  1  1  7 */ assign n330 = n331;

endmodule

