// Reading file 'blink.asc'..

module chip (input io_0_8_1, output io_13_6_1);

wire io_0_8_1;
// (0, 0, 'glb_netwk_6')
// (0, 5, 'span4_vert_t_14')
// (0, 6, 'span4_vert_b_14')
// (0, 7, 'span4_vert_b_10')
// (0, 8, 'fabout')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'local_g1_6')
// (0, 8, 'span4_vert_b_6')
// (0, 9, 'span4_vert_b_2')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (11, 3, 'lutff_global/clk')
// (12, 3, 'lutff_global/clk')
// (12, 4, 'lutff_global/clk')
// (12, 5, 'lutff_global/clk')

reg n2 = 0;
// (10, 2, 'neigh_op_tnr_3')
// (10, 3, 'neigh_op_rgt_3')
// (10, 4, 'neigh_op_bnr_3')
// (11, 2, 'neigh_op_top_3')
// (11, 3, 'local_g0_3')
// (11, 3, 'lutff_3/in_0')
// (11, 3, 'lutff_3/out')
// (11, 4, 'neigh_op_bot_3')
// (12, 2, 'neigh_op_tnl_3')
// (12, 3, 'local_g1_3')
// (12, 3, 'lutff_0/in_2')
// (12, 3, 'lutff_1/in_3')
// (12, 3, 'neigh_op_lft_3')
// (12, 4, 'neigh_op_bnl_3')

reg n3 = 0;
// (11, 2, 'neigh_op_tnr_1')
// (11, 3, 'neigh_op_rgt_1')
// (11, 4, 'neigh_op_bnr_1')
// (12, 2, 'neigh_op_top_1')
// (12, 3, 'local_g2_1')
// (12, 3, 'lutff_1/in_2')
// (12, 3, 'lutff_1/out')
// (12, 4, 'neigh_op_bot_1')
// (13, 2, 'logic_op_tnl_1')
// (13, 3, 'logic_op_lft_1')
// (13, 4, 'logic_op_bnl_1')

reg n4 = 0;
// (11, 2, 'neigh_op_tnr_2')
// (11, 3, 'neigh_op_rgt_2')
// (11, 4, 'neigh_op_bnr_2')
// (12, 2, 'neigh_op_top_2')
// (12, 3, 'local_g1_2')
// (12, 3, 'lutff_2/in_1')
// (12, 3, 'lutff_2/out')
// (12, 4, 'neigh_op_bot_2')
// (13, 2, 'logic_op_tnl_2')
// (13, 3, 'logic_op_lft_2')
// (13, 4, 'logic_op_bnl_2')

reg n5 = 0;
// (11, 2, 'neigh_op_tnr_3')
// (11, 3, 'neigh_op_rgt_3')
// (11, 4, 'neigh_op_bnr_3')
// (12, 2, 'neigh_op_top_3')
// (12, 3, 'local_g0_3')
// (12, 3, 'lutff_3/in_2')
// (12, 3, 'lutff_3/out')
// (12, 4, 'neigh_op_bot_3')
// (13, 2, 'logic_op_tnl_3')
// (13, 3, 'logic_op_lft_3')
// (13, 4, 'logic_op_bnl_3')

reg n6 = 0;
// (11, 2, 'neigh_op_tnr_4')
// (11, 3, 'neigh_op_rgt_4')
// (11, 4, 'neigh_op_bnr_4')
// (12, 2, 'neigh_op_top_4')
// (12, 3, 'local_g3_4')
// (12, 3, 'lutff_4/in_1')
// (12, 3, 'lutff_4/out')
// (12, 4, 'neigh_op_bot_4')
// (13, 2, 'logic_op_tnl_4')
// (13, 3, 'logic_op_lft_4')
// (13, 4, 'logic_op_bnl_4')

reg n7 = 0;
// (11, 2, 'neigh_op_tnr_5')
// (11, 3, 'neigh_op_rgt_5')
// (11, 4, 'neigh_op_bnr_5')
// (12, 2, 'neigh_op_top_5')
// (12, 3, 'local_g2_5')
// (12, 3, 'lutff_5/in_2')
// (12, 3, 'lutff_5/out')
// (12, 4, 'neigh_op_bot_5')
// (13, 2, 'logic_op_tnl_5')
// (13, 3, 'logic_op_lft_5')
// (13, 4, 'logic_op_bnl_5')

reg n8 = 0;
// (11, 2, 'neigh_op_tnr_6')
// (11, 3, 'neigh_op_rgt_6')
// (11, 4, 'neigh_op_bnr_6')
// (12, 2, 'neigh_op_top_6')
// (12, 3, 'local_g0_6')
// (12, 3, 'lutff_6/in_2')
// (12, 3, 'lutff_6/out')
// (12, 4, 'neigh_op_bot_6')
// (13, 2, 'logic_op_tnl_6')
// (13, 3, 'logic_op_lft_6')
// (13, 4, 'logic_op_bnl_6')

reg n9 = 0;
// (11, 2, 'neigh_op_tnr_7')
// (11, 3, 'neigh_op_rgt_7')
// (11, 4, 'neigh_op_bnr_7')
// (12, 2, 'neigh_op_top_7')
// (12, 3, 'local_g2_7')
// (12, 3, 'lutff_7/in_2')
// (12, 3, 'lutff_7/out')
// (12, 4, 'neigh_op_bot_7')
// (13, 2, 'logic_op_tnl_7')
// (13, 3, 'logic_op_lft_7')
// (13, 4, 'logic_op_bnl_7')

reg n10 = 0;
// (11, 3, 'neigh_op_tnr_0')
// (11, 4, 'neigh_op_rgt_0')
// (11, 5, 'neigh_op_bnr_0')
// (12, 3, 'neigh_op_top_0')
// (12, 4, 'local_g3_0')
// (12, 4, 'lutff_0/in_1')
// (12, 4, 'lutff_0/out')
// (12, 5, 'neigh_op_bot_0')
// (13, 3, 'logic_op_tnl_0')
// (13, 4, 'logic_op_lft_0')
// (13, 5, 'logic_op_bnl_0')

reg n11 = 0;
// (11, 3, 'neigh_op_tnr_1')
// (11, 4, 'neigh_op_rgt_1')
// (11, 5, 'neigh_op_bnr_1')
// (12, 3, 'neigh_op_top_1')
// (12, 4, 'local_g3_1')
// (12, 4, 'lutff_1/in_1')
// (12, 4, 'lutff_1/out')
// (12, 5, 'neigh_op_bot_1')
// (13, 3, 'logic_op_tnl_1')
// (13, 4, 'logic_op_lft_1')
// (13, 5, 'logic_op_bnl_1')

reg n12 = 0;
// (11, 3, 'neigh_op_tnr_2')
// (11, 4, 'neigh_op_rgt_2')
// (11, 5, 'neigh_op_bnr_2')
// (12, 3, 'neigh_op_top_2')
// (12, 4, 'local_g3_2')
// (12, 4, 'lutff_2/in_1')
// (12, 4, 'lutff_2/out')
// (12, 5, 'neigh_op_bot_2')
// (13, 3, 'logic_op_tnl_2')
// (13, 4, 'logic_op_lft_2')
// (13, 5, 'logic_op_bnl_2')

reg n13 = 0;
// (11, 3, 'neigh_op_tnr_3')
// (11, 4, 'neigh_op_rgt_3')
// (11, 5, 'neigh_op_bnr_3')
// (12, 3, 'neigh_op_top_3')
// (12, 4, 'local_g2_3')
// (12, 4, 'lutff_3/in_2')
// (12, 4, 'lutff_3/out')
// (12, 5, 'neigh_op_bot_3')
// (13, 3, 'logic_op_tnl_3')
// (13, 4, 'logic_op_lft_3')
// (13, 5, 'logic_op_bnl_3')

reg n14 = 0;
// (11, 3, 'neigh_op_tnr_4')
// (11, 4, 'neigh_op_rgt_4')
// (11, 5, 'neigh_op_bnr_4')
// (12, 3, 'neigh_op_top_4')
// (12, 4, 'local_g2_4')
// (12, 4, 'lutff_4/in_2')
// (12, 4, 'lutff_4/out')
// (12, 5, 'neigh_op_bot_4')
// (13, 3, 'logic_op_tnl_4')
// (13, 4, 'logic_op_lft_4')
// (13, 5, 'logic_op_bnl_4')

reg n15 = 0;
// (11, 3, 'neigh_op_tnr_5')
// (11, 4, 'neigh_op_rgt_5')
// (11, 5, 'neigh_op_bnr_5')
// (12, 3, 'neigh_op_top_5')
// (12, 4, 'local_g0_5')
// (12, 4, 'lutff_5/in_2')
// (12, 4, 'lutff_5/out')
// (12, 5, 'neigh_op_bot_5')
// (13, 3, 'logic_op_tnl_5')
// (13, 4, 'logic_op_lft_5')
// (13, 5, 'logic_op_bnl_5')

reg n16 = 0;
// (11, 3, 'neigh_op_tnr_6')
// (11, 4, 'neigh_op_rgt_6')
// (11, 5, 'neigh_op_bnr_6')
// (12, 3, 'neigh_op_top_6')
// (12, 4, 'local_g3_6')
// (12, 4, 'lutff_6/in_1')
// (12, 4, 'lutff_6/out')
// (12, 5, 'neigh_op_bot_6')
// (13, 3, 'logic_op_tnl_6')
// (13, 4, 'logic_op_lft_6')
// (13, 5, 'logic_op_bnl_6')

reg n17 = 0;
// (11, 3, 'neigh_op_tnr_7')
// (11, 4, 'neigh_op_rgt_7')
// (11, 5, 'neigh_op_bnr_7')
// (12, 3, 'neigh_op_top_7')
// (12, 4, 'local_g0_7')
// (12, 4, 'lutff_7/in_2')
// (12, 4, 'lutff_7/out')
// (12, 5, 'neigh_op_bot_7')
// (13, 3, 'logic_op_tnl_7')
// (13, 4, 'logic_op_lft_7')
// (13, 5, 'logic_op_bnl_7')

reg n18 = 0;
// (11, 4, 'neigh_op_tnr_0')
// (11, 5, 'neigh_op_rgt_0')
// (11, 6, 'neigh_op_bnr_0')
// (12, 4, 'neigh_op_top_0')
// (12, 5, 'local_g0_0')
// (12, 5, 'lutff_0/in_2')
// (12, 5, 'lutff_0/out')
// (12, 6, 'neigh_op_bot_0')
// (13, 4, 'logic_op_tnl_0')
// (13, 5, 'logic_op_lft_0')
// (13, 6, 'logic_op_bnl_0')

reg n19 = 0;
// (11, 4, 'neigh_op_tnr_1')
// (11, 5, 'neigh_op_rgt_1')
// (11, 6, 'neigh_op_bnr_1')
// (12, 4, 'neigh_op_top_1')
// (12, 5, 'local_g2_1')
// (12, 5, 'lutff_1/in_2')
// (12, 5, 'lutff_1/out')
// (12, 6, 'neigh_op_bot_1')
// (13, 4, 'logic_op_tnl_1')
// (13, 5, 'logic_op_lft_1')
// (13, 6, 'logic_op_bnl_1')

reg n20 = 0;
// (11, 4, 'neigh_op_tnr_2')
// (11, 5, 'neigh_op_rgt_2')
// (11, 6, 'neigh_op_bnr_2')
// (12, 4, 'neigh_op_top_2')
// (12, 5, 'local_g0_2')
// (12, 5, 'lutff_2/in_2')
// (12, 5, 'lutff_2/out')
// (12, 6, 'neigh_op_bot_2')
// (13, 4, 'logic_op_tnl_2')
// (13, 5, 'logic_op_lft_2')
// (13, 6, 'logic_op_bnl_2')

reg n21 = 0;
// (11, 4, 'neigh_op_tnr_3')
// (11, 5, 'neigh_op_rgt_3')
// (11, 6, 'neigh_op_bnr_3')
// (12, 4, 'neigh_op_top_3')
// (12, 5, 'local_g0_3')
// (12, 5, 'lutff_3/in_2')
// (12, 5, 'lutff_3/out')
// (12, 6, 'neigh_op_bot_3')
// (13, 4, 'logic_op_tnl_3')
// (13, 5, 'logic_op_lft_3')
// (13, 6, 'logic_op_bnl_3')

reg n22 = 0;
// (11, 4, 'neigh_op_tnr_4')
// (11, 5, 'neigh_op_rgt_4')
// (11, 6, 'neigh_op_bnr_4')
// (12, 4, 'neigh_op_top_4')
// (12, 5, 'local_g0_4')
// (12, 5, 'lutff_4/in_2')
// (12, 5, 'lutff_4/out')
// (12, 6, 'neigh_op_bot_4')
// (13, 4, 'logic_op_tnl_4')
// (13, 5, 'logic_op_lft_4')
// (13, 6, 'logic_op_bnl_4')

reg n23 = 0;
// (11, 4, 'neigh_op_tnr_5')
// (11, 5, 'neigh_op_rgt_5')
// (11, 6, 'neigh_op_bnr_5')
// (12, 4, 'neigh_op_top_5')
// (12, 5, 'local_g0_5')
// (12, 5, 'lutff_5/in_2')
// (12, 5, 'lutff_5/out')
// (12, 6, 'neigh_op_bot_5')
// (13, 4, 'logic_op_tnl_5')
// (13, 5, 'logic_op_lft_5')
// (13, 6, 'logic_op_bnl_5')

reg n24 = 0;
// (11, 4, 'neigh_op_tnr_6')
// (11, 5, 'neigh_op_rgt_6')
// (11, 6, 'neigh_op_bnr_6')
// (12, 4, 'neigh_op_top_6')
// (12, 5, 'local_g2_6')
// (12, 5, 'lutff_6/in_2')
// (12, 5, 'lutff_6/out')
// (12, 6, 'neigh_op_bot_6')
// (13, 4, 'logic_op_tnl_6')
// (13, 5, 'logic_op_lft_6')
// (13, 6, 'logic_op_bnl_6')

reg io_13_6_1 = 0;
// (11, 4, 'neigh_op_tnr_7')
// (11, 5, 'neigh_op_rgt_7')
// (11, 6, 'neigh_op_bnr_7')
// (12, 4, 'neigh_op_top_7')
// (12, 5, 'local_g0_7')
// (12, 5, 'lutff_7/in_2')
// (12, 5, 'lutff_7/out')
// (12, 6, 'neigh_op_bot_7')
// (13, 4, 'logic_op_tnl_7')
// (13, 5, 'logic_op_lft_7')
// (13, 6, 'io_1/D_OUT_0')
// (13, 6, 'io_1/PAD')
// (13, 6, 'local_g0_7')
// (13, 6, 'logic_op_bnl_7')

wire n26;
// (12, 3, 'lutff_1/cout')
// (12, 3, 'lutff_2/in_3')

wire n27;
// (12, 3, 'lutff_2/cout')
// (12, 3, 'lutff_3/in_3')

wire n28;
// (12, 3, 'lutff_3/cout')
// (12, 3, 'lutff_4/in_3')

wire n29;
// (12, 3, 'lutff_4/cout')
// (12, 3, 'lutff_5/in_3')

wire n30;
// (12, 3, 'lutff_5/cout')
// (12, 3, 'lutff_6/in_3')

wire n31;
// (12, 3, 'lutff_6/cout')
// (12, 3, 'lutff_7/in_3')

wire n32;
// (12, 3, 'lutff_7/cout')
// (12, 4, 'carry_in')
// (12, 4, 'carry_in_mux')
// (12, 4, 'lutff_0/in_3')

wire n33;
// (12, 4, 'lutff_0/cout')
// (12, 4, 'lutff_1/in_3')

wire n34;
// (12, 4, 'lutff_1/cout')
// (12, 4, 'lutff_2/in_3')

wire n35;
// (12, 4, 'lutff_2/cout')
// (12, 4, 'lutff_3/in_3')

wire n36;
// (12, 4, 'lutff_3/cout')
// (12, 4, 'lutff_4/in_3')

wire n37;
// (12, 4, 'lutff_4/cout')
// (12, 4, 'lutff_5/in_3')

wire n38;
// (12, 4, 'lutff_5/cout')
// (12, 4, 'lutff_6/in_3')

wire n39;
// (12, 4, 'lutff_6/cout')
// (12, 4, 'lutff_7/in_3')

wire n40;
// (12, 4, 'lutff_7/cout')
// (12, 5, 'carry_in')
// (12, 5, 'carry_in_mux')
// (12, 5, 'lutff_0/in_3')

wire n41;
// (12, 5, 'lutff_0/cout')
// (12, 5, 'lutff_1/in_3')

wire n42;
// (12, 5, 'lutff_1/cout')
// (12, 5, 'lutff_2/in_3')

wire n43;
// (12, 5, 'lutff_2/cout')
// (12, 5, 'lutff_3/in_3')

wire n44;
// (12, 5, 'lutff_3/cout')
// (12, 5, 'lutff_4/in_3')

wire n45;
// (12, 5, 'lutff_4/cout')
// (12, 5, 'lutff_5/in_3')

wire n46;
// (12, 5, 'lutff_5/cout')
// (12, 5, 'lutff_6/in_3')

wire n47;
// (12, 5, 'lutff_6/cout')
// (12, 5, 'lutff_7/in_3')

wire n48;
// (12, 3, 'lutff_0/cout')

wire n49;
// (12, 4, 'lutff_2/lout')

wire n50;
// (12, 4, 'lutff_5/lout')

wire n51;
// (12, 3, 'lutff_0/out')

wire n52;
// (12, 3, 'lutff_0/lout')

wire n53;
// (12, 3, 'carry_in_mux')

// Carry-In for (12 3)
assign n53 = 1;

wire n54;
// (12, 3, 'lutff_3/lout')

wire n55;
// (12, 5, 'lutff_0/lout')

wire n56;
// (12, 3, 'lutff_6/lout')

wire n57;
// (12, 5, 'lutff_3/lout')

wire n58;
// (12, 5, 'lutff_6/lout')

wire n59;
// (12, 4, 'lutff_1/lout')

wire n60;
// (12, 4, 'lutff_7/lout')

wire n61;
// (12, 4, 'lutff_4/lout')

wire n62;
// (11, 3, 'lutff_3/lout')

wire n63;
// (12, 3, 'lutff_5/lout')

wire n64;
// (12, 5, 'lutff_2/lout')

wire n65;
// (12, 3, 'lutff_2/lout')

wire n66;
// (12, 5, 'lutff_5/lout')

wire n67;
// (12, 4, 'lutff_0/lout')

wire n68;
// (12, 4, 'lutff_3/lout')

wire n69;
// (12, 4, 'lutff_6/lout')

wire n70;
// (12, 3, 'lutff_1/lout')

wire n71;
// (12, 3, 'lutff_7/lout')

wire n72;
// (12, 3, 'lutff_4/lout')

wire n73;
// (12, 5, 'lutff_1/lout')

wire n74;
// (12, 5, 'lutff_7/lout')

wire n75;
// (12, 5, 'lutff_4/lout')

assign n52 = /* LUT   12  3  0 */ 1'b0;
assign n49 = /* LUT   12  4  2 */ (n34 ? !n12 : n12);
assign n50 = /* LUT   12  4  5 */ (n37 ? !n15 : n15);
assign n54 = /* LUT   12  3  3 */ (n27 ? !n5 : n5);
assign n55 = /* LUT   12  5  0 */ (n40 ? !n18 : n18);
assign n56 = /* LUT   12  3  6 */ (n30 ? !n8 : n8);
assign n57 = /* LUT   12  5  3 */ (n43 ? !n21 : n21);
assign n58 = /* LUT   12  5  6 */ (n46 ? !n24 : n24);
assign n59 = /* LUT   12  4  1 */ (n33 ? !n11 : n11);
assign n60 = /* LUT   12  4  7 */ (n39 ? !n17 : n17);
assign n61 = /* LUT   12  4  4 */ (n36 ? !n14 : n14);
assign n62 = /* LUT   11  3  3 */ !n2;
assign n63 = /* LUT   12  3  5 */ (n29 ? !n7 : n7);
assign n64 = /* LUT   12  5  2 */ (n42 ? !n20 : n20);
assign n65 = /* LUT   12  3  2 */ (n26 ? !n4 : n4);
assign n66 = /* LUT   12  5  5 */ (n45 ? !n23 : n23);
assign n67 = /* LUT   12  4  0 */ (n32 ? !n10 : n10);
assign n68 = /* LUT   12  4  3 */ (n35 ? !n13 : n13);
assign n69 = /* LUT   12  4  6 */ (n38 ? !n16 : n16);
assign n70 = /* LUT   12  3  1 */ (n2 ? !n3 : n3);
assign n71 = /* LUT   12  3  7 */ (n31 ? !n9 : n9);
assign n72 = /* LUT   12  3  4 */ (n28 ? !n6 : n6);
assign n73 = /* LUT   12  5  1 */ (n41 ? !n19 : n19);
assign n74 = /* LUT   12  5  7 */ (n47 ? !io_13_6_1 : io_13_6_1);
assign n75 = /* LUT   12  5  4 */ (n44 ? !n22 : n22);
assign n35 = /* CARRY 12  4  2 */ (n12 & 1'b0) | ((n12 | 1'b0) & n34);
assign n38 = /* CARRY 12  4  5 */ (1'b0 & n15) | ((1'b0 | n15) & n37);
assign n48 = /* CARRY 12  3  0 */ (1'b0 & n2) | ((1'b0 | n2) & n53);
assign n28 = /* CARRY 12  3  3 */ (1'b0 & n5) | ((1'b0 | n5) & n27);
assign n41 = /* CARRY 12  5  0 */ (1'b0 & n18) | ((1'b0 | n18) & n40);
assign n31 = /* CARRY 12  3  6 */ (1'b0 & n8) | ((1'b0 | n8) & n30);
assign n44 = /* CARRY 12  5  3 */ (1'b0 & n21) | ((1'b0 | n21) & n43);
assign n47 = /* CARRY 12  5  6 */ (1'b0 & n24) | ((1'b0 | n24) & n46);
assign n34 = /* CARRY 12  4  1 */ (n11 & 1'b0) | ((n11 | 1'b0) & n33);
assign n40 = /* CARRY 12  4  7 */ (1'b0 & n17) | ((1'b0 | n17) & n39);
assign n37 = /* CARRY 12  4  4 */ (1'b0 & n14) | ((1'b0 | n14) & n36);
assign n30 = /* CARRY 12  3  5 */ (1'b0 & n7) | ((1'b0 | n7) & n29);
assign n43 = /* CARRY 12  5  2 */ (1'b0 & n20) | ((1'b0 | n20) & n42);
assign n27 = /* CARRY 12  3  2 */ (n4 & 1'b0) | ((n4 | 1'b0) & n26);
assign n46 = /* CARRY 12  5  5 */ (1'b0 & n23) | ((1'b0 | n23) & n45);
assign n33 = /* CARRY 12  4  0 */ (n10 & 1'b0) | ((n10 | 1'b0) & n32);
assign n36 = /* CARRY 12  4  3 */ (1'b0 & n13) | ((1'b0 | n13) & n35);
assign n39 = /* CARRY 12  4  6 */ (n16 & 1'b0) | ((n16 | 1'b0) & n38);
assign n26 = /* CARRY 12  3  1 */ (1'b0 & n3) | ((1'b0 | n3) & n48);
assign n32 = /* CARRY 12  3  7 */ (1'b0 & n9) | ((1'b0 | n9) & n31);
assign n29 = /* CARRY 12  3  4 */ (n6 & 1'b0) | ((n6 | 1'b0) & n28);
assign n42 = /* CARRY 12  5  1 */ (1'b0 & n19) | ((1'b0 | n19) & n41);
assign n45 = /* CARRY 12  5  4 */ (1'b0 & n22) | ((1'b0 | n22) & n44);
/* FF 12  4  2 */ always @(posedge io_0_8_1) if (1'b1) n12 <= 1'b0 ? 1'b0 : n49;
/* FF 12  4  5 */ always @(posedge io_0_8_1) if (1'b1) n15 <= 1'b0 ? 1'b0 : n50;
/* FF 12  3  0 */ assign n51 = n52;
/* FF 12  3  3 */ always @(posedge io_0_8_1) if (1'b1) n5 <= 1'b0 ? 1'b0 : n54;
/* FF 12  5  0 */ always @(posedge io_0_8_1) if (1'b1) n18 <= 1'b0 ? 1'b0 : n55;
/* FF 12  3  6 */ always @(posedge io_0_8_1) if (1'b1) n8 <= 1'b0 ? 1'b0 : n56;
/* FF 12  5  3 */ always @(posedge io_0_8_1) if (1'b1) n21 <= 1'b0 ? 1'b0 : n57;
/* FF 12  5  6 */ always @(posedge io_0_8_1) if (1'b1) n24 <= 1'b0 ? 1'b0 : n58;
/* FF 12  4  1 */ always @(posedge io_0_8_1) if (1'b1) n11 <= 1'b0 ? 1'b0 : n59;
/* FF 12  4  7 */ always @(posedge io_0_8_1) if (1'b1) n17 <= 1'b0 ? 1'b0 : n60;
/* FF 12  4  4 */ always @(posedge io_0_8_1) if (1'b1) n14 <= 1'b0 ? 1'b0 : n61;
/* FF 11  3  3 */ always @(posedge io_0_8_1) if (1'b1) n2 <= 1'b0 ? 1'b0 : n62;
/* FF 12  3  5 */ always @(posedge io_0_8_1) if (1'b1) n7 <= 1'b0 ? 1'b0 : n63;
/* FF 12  5  2 */ always @(posedge io_0_8_1) if (1'b1) n20 <= 1'b0 ? 1'b0 : n64;
/* FF 12  3  2 */ always @(posedge io_0_8_1) if (1'b1) n4 <= 1'b0 ? 1'b0 : n65;
/* FF 12  5  5 */ always @(posedge io_0_8_1) if (1'b1) n23 <= 1'b0 ? 1'b0 : n66;
/* FF 12  4  0 */ always @(posedge io_0_8_1) if (1'b1) n10 <= 1'b0 ? 1'b0 : n67;
/* FF 12  4  3 */ always @(posedge io_0_8_1) if (1'b1) n13 <= 1'b0 ? 1'b0 : n68;
/* FF 12  4  6 */ always @(posedge io_0_8_1) if (1'b1) n16 <= 1'b0 ? 1'b0 : n69;
/* FF 12  3  1 */ always @(posedge io_0_8_1) if (1'b1) n3 <= 1'b0 ? 1'b0 : n70;
/* FF 12  3  7 */ always @(posedge io_0_8_1) if (1'b1) n9 <= 1'b0 ? 1'b0 : n71;
/* FF 12  3  4 */ always @(posedge io_0_8_1) if (1'b1) n6 <= 1'b0 ? 1'b0 : n72;
/* FF 12  5  1 */ always @(posedge io_0_8_1) if (1'b1) n19 <= 1'b0 ? 1'b0 : n73;
/* FF 12  5  7 */ always @(posedge io_0_8_1) if (1'b1) io_13_6_1 <= 1'b0 ? 1'b0 : n74;
/* FF 12  5  4 */ always @(posedge io_0_8_1) if (1'b1) n22 <= 1'b0 ? 1'b0 : n75;

endmodule

